PK   ��X)$�  �     cirkitFile.json�][�㸱�+�%,G�S���Mp�f���a�ѠDj['nˑ幜���C�wI��.v� �Ơ���E�cU�TR�4�Y<ucޛfUՋ�-b�ɣj�u|5�N��⡭~k��qr��}O�OK��Ӳ^�E���*E
�	�'���J�$5�(�a9C�!�ܾ��>���1���ةec6��,3:A8g	�M�(�e�4S)����̣�L1��yB�D����S��ʼ�ER;� �Dk�A���Kn���	��H(!"ɸ�	.�+��Al��gИ����Ɛ�3ஆZ�Y@@����Q ?�s � �K ?�?uK@�a �0�3!��� �bw�h�a����ń���a��8p�b�n���J����wk�짞u<M��&�
m�,Cy"�.���]rRpoh�}�4�g��
�@=�,[`���g��!󉄳'Th��kC%2H�������A �[� v�a	b�ە���+�~�5[�B|0�o��n�7h����0n�x����<���Yxz̂��+�d���<�z��(3̏ �c�}'�g�lw��}�70���E&�_�ޢ��0�;�C���qB���(RH)�I)K�EE��2"�`�q��,�"�7zQ��8�E4��8Fq �D12��8(�qP�#��8(�qP�is�;2701[�,!b��A1��b��"�C�~��K34A���)4�aD,���.!4�A�ŭ�ъ��H�E�Lgp����:�7��	�ڰ8�\�phv'����*4�A�E#����3�R`�����f���=��r��Z�h&`a�m���L \
�"�D�B�HaQ��(RD)2��,�"�7zQ��8�Eq �� Ł0��a�(�q�H68�q�8(�qP���A1��b�$��Eg�R��rqCg�R.n��L \����	�K����3P	�q�{9�	�D�����L�Y1�� �����	�K����H$4 �rqD�� ��c]�L�Ǐ�"��'��O'�Ƭ�sU�P-�F�fr�n���Li�J�%)�1��<SIV�bE�N�	ר<�g�CU�u9��yP�
��S4^3��=�f���3�!��!c��;�]A2Y���
�!={f;���ol���:3P ���0�����a�$�ك��JR��:���gX��س������|���ȸ1O�{�����Y-�Zs�:) ���*�:�s��s�at�Bt!�9P	P���nF���\�!���BzV�����P��p; �;�g�o_}|u_���  ��/�BO�gx�*P#p	�pP�+ </�U�5��p��g�6�#� >K�Ӵj��Z��P���]���Q]WZ�� �M��c ?�[���g�KR{�<h�M퉃q��5�Z�'� +�`,C���hFP8w% *�C� 	 E"�"��*��D<bY�YÁ<`
p �K�P�b(l1�
[r����=w�g�O�BFG����rӞ8H�9��2`jO�'K\�
��3�+���.8	�8��ᥧa�4�5̞����o� ���9���=}<�.�B�'������y�Kp�jO$]7�]��=i[\��籤�u�=�x�\���=�zSi�X��W.���ݻ��8��Qr�m.��6�nF�4t.�Aw����1r�ȑ#G�r�q�N����;�.���Z����;�8H�
ѐ�U}�gȆ=�iB@��e
��I/!�8b��Xo��0�C��捋=h�^��JE�C{&ȣ�w��	�zM�7�%0c�Za9�=��QB� ��ɡO��r��Ua�7�/w�
3�����:�a$z�5�ptǀ^��%�-�����K�!���{fOݺǕ�*7s�{������m�^�6�a�6�a�6�a�6�a�6�aS�mJ�Mb�$�Mr�$�Mٶ)4�]_h����X��yc��kոZֲ~�W�v�[���A��^��]z��KӴ��������V�v�j�j�Uh���w�:��W����n�ܼ���db?��?-��r'�����m\���jU�s��֘�����m۬�ԓZ�KU���4�8&;�ds+2�&�m;��j�?����t���	f�ϩ���و_猦$����i��ۍ�{E0A���~���1��ĞbZ�(6���2�I�TV���4i��['�j���.�;,ŌM1O炙�N���,�� j�B��^*�NZ𡅥����|-��Q��^��C�n�R~����39�Ύ�����zv�N��:�|0���<:���E��16Ǜ��9޶���ed��-#s�m�qg��ۯ��iYϵi��ﺽ}7�����e���n2��T��B�!D3���n�e��'J�BD�yGo>.�5
��>��lx3AT���N�	��'k� �1s;q������a*N04���D��&e��,�9��Y,��q�y��6Ltf�+W�$G&�>����Y�0�p�f�q"~�sr��G��|�X���d���sT$,͕��)K0�B�2/RJO��{�4u���,�'MIP�'\b��S�&����X��H!؈�����kS����Z�Tq;���@�I�s�u�S��v���Tm�3��ڶr�;����|�I�^�U����	��C�q�ۺi��ucV�mۗ)r@���܌�kVmEo�I)n�xY��Z5)�8��ӒS;S���	ĕ18���[K�Ki�pILf�*Y10��r@H�yB�ȓQf��B�IԢ�^�)c�RA�Ć�VaTdIn\hktZ2Α΋� +6_�&��J߬L�^��O7���77�����S�n6-7����4fz��7�zqS[�uk��/��:A���ň��,�j��:���37E�A����4�N6���.�|{�F3L�������W��ҮuU�=��ȌX�@cD��W|�*�u�޼Y��#� Y|�O9�3;�4C'���9�	NI�!���$�2���((S��������v���(�(l�d����]��{�B(�e�X�i³�W�m�c��S��4+�T�yb2LF�L���D3a�
�C��}����XM]�ҋ�Rb�c[,�,���0#d��Q4	<�"z��_ EA7!P$p"k��� ;�4�8x~��M��3�����~����:F���&S��	��V��W�Bq!�ۺ)�3�P^j�IA1e���;y!��Č�b���'��ѐ��YJr{��:I��:�L�[b{�%3�q���:2�f�Y��Βe��ow�Y2�R{��g�Y��F 	�oH� �;Y���Y�	+��f��9���p{HJ������sJ�n�����%�Q{��u�tg_���`+�`Fw�R�v���~����$�k=J�7�`q�Ln�1r���D/] vN���tϱ;}��͸��ՃY "�ѓ��n
#�y��ۋjЩB��fj+�>����t7:�ѧ�d�L�1����H�m�H<t���ܞ��.:��4�.e[����mm�$A�Yk�e���]��m�]$����,p8��9�Gӥo'C�ԞB��x���T�+�Pţ���S�oӶ�~�̇�W'�{�݁ў|���]��)ͮPӾ��s���o��}VV���NV�>�U9+��[�բ}���N�=0�M\����k��s�+w����ݥ���z8�:���u0],��`ؖ��������o�C�eg��^vw�q�e?I�t��T�!�N��e�/��6̻���E�T����S�Bh�X�B�G��!B$����E��
���eg�����\�gP�Ƶ�ݑ�^A�NJD�!(��/2���s�vW§�3~6��]^�Z*F� {�%�n�vq��g9����Q[��3��(.8}� <�!�Ů��g�"ڞ�j�  ^��@�B�  ^�ݕ@<M��I���K�_��_[�i{"&6b�t�5�u��/Ӹ-�ܺ��������T7�a>�����
�@�s�
��ٞ+�x�j�lϳ���C����@�Z�G�uc�TE�P�Y��2��JO�F�BCݫ�aO����2�.�Qw�|�.?�Y���T��q>�����i�E��]�Z��?/�D'a����SnS��ÝlY���R�E�&�Z�E�I�d˻�T������",z��a���~�j�R��Y�C�ՙ5��g�S��Ķ�"���g�����+T����JVv�v�L{��Q��_��f�]�F5��T��Z�Tj���:��/����Z������Mk�����P�M���h0������ɗ�PK   
��X[�o��� �� /   images/055d5e06-61e9-48ec-9da3-6ebf1aca914f.png�{�S�-4@�܃-��H����{��	�I���N�w��܂�./<��������jj���z���{�9=��T��S>GAA�WT��@AA=�wbc>���G<]p��\QP޾�w�zJx����(�Hize =v��ၰ�uŤR�e?��å��A�A2r�Φ�]��TQX�V�Üc^b�T�mx���܌��б7�����^�:�OqD�w���Zo���Q]����J�سD�ms��mj�?������X�Es)5����Z��Su�(�?n���?\J<G���<����CqS;O�M�)�
��?�M�H���"�ү�t�����	�GϞI<T>b{?�H�o$���B=��_���MB�Ћ�z%���M��Vz��p���
TO@/&��� ����``ʽb��2�Qa��IZ<=f��b���O=����k�M����� P�q��iW����r}�<&E����(��]y!1�5a�-HabJ$"i`��)�l�EJa�|e�3����3�NT�F�?��[8��?��L@�S�����|��6���I�_��:o�a3Dޕc�uL�$g	��6n$�51���g��٦�+�\>� �(���L�,��o�S"-�!��@J
 ��6����ߺv�%%�3�졹Y�*<�%��E�Y���"���"V5�C�/�D5�{��Ձޥ\F�P�����n~����'j��UH�8�˪�Z���`t���j�F��:_�ݹ�ø��=F}
5i�\�{lIX�aq��r�����S�&A�����8 ���u�b"i6:4/묫PST\]D��vQ1W��I��@�b��eu�gF�q�@*2C��v�U�:O�n�EL��,ٸ��#�n���1����}3ڝ49e�@�}̗û�ӠRȯ
N��>r�I\��sS��լ�l��K:va�s�լ�b�(l���E����ɜ\��-���q��_�b�Ӷؔ�Q�^Yx/?����}>���B���\K���^e�;���?y@G���:�|���Ni�_g�_G�W*�_�;X�@���$�Ӏ�	b�?�a��}��{)�)E�n$o���ê���?��8�g`���v�K���U�"jc�$�黑�Fu�ˋ��wJ��v�R-l��"��_�i�Eە��7� �s�UY;?���%��"�j:��Af"=³�112-A�	�����M�>&�"p��d݌�o��#�ŝ����Ú�x��]�	��$�no��虯�^g1�_�I2H)O�)��)������/�]���j��I�LS��Y�@J� ��)���4��&`���v:���i~Zӳ5�C��e��9ˇ4�x�4��k3�O9��/G�0�7�?��!���,��jiaO!Mіk_M��wx/~ ��%� ��_d�.��c��J�A$`JT�o�a[�A�>�L��'�%h�]��L~��;�w���"z��H�Q��3&��0"ybCgf�t��lZjC��S�E��������p��g}�ONN9TB��0����յ����=%��I^!�M��"�1a�a Ǘ�#��J&�[=���|�\�dh���psp1��.�v��"��@�i����1�.�N0���H��P�,I����2J$-���"JV��`����>�����Z
T)������7پ���|�9󦖮I��n�^DF\Щ+�Kh�>����(;�p�.�"�� q�C��|6{�Lb�����n����|�&���d�qE����0ֱ�>H�#�+����ʨ�������C��9f�]Λ�P���K����]�|)���[c����^f�}3�3�e��-?���+�fQ��+V����N��!��lG�
��V���x��l~J)�q�	����H�����oG��:K�[j𐨜N�pN���V!�{[���w
�ґye�^���b����ؕ��I���ၾ���2����3p6?�I�씓U#]l���k���J�x�u��4l��u�r�<l�>"�>�"mF�%��ؿ�C�qm/̄�o{4����R�ZHrD�0�Y"�CC	Q�ٻÿ5��R�ɰ�H)�ZГ;����.��
<�B����o��4���=�w�ϫ���STy����$�#ڰ��R�.���<Y5٪�{&6e�E�E��5"i5��ce6��^Kx�����#���ur���L��x�p�~ą�OR��ƪ���{@��J:�DaB�ǽJ׳F��V�_�V�����11�%�A2
��?ɤ�j1U.�M,I�߂\	��Xܣ4�W�Y#^���`�`���@�����]$�r��Ɓ�Z|��?�X3%\c^*E�\�4��E��U�FG���8��m|�>�8:������PK��A���*y�r,�\W�W%A[����^�����0� ��t���8b6Ӏ����W�$�P$�k%����df���󑄐��ȲΓ��6���⹇�;��FX�H��:��-�f���oD3����/ͪ�5�/1!�
<
�d�
/|����mQ|��w��/بgk)>�uR�/�賧�M:@������hNhU>1��cC7��ⵘq��"7�¤��joV��:�!}��n�vv��z��骁E��B�tc%4$�	8�XX�џ���s$`��j��w<<P���=���>��F�"��mp�j��!�_9d�a$��Jv$)�J�c�]��p�G��ݘ���exr ���*\"�J��ε��t^Cd,ϔaw����)�>U%��Ώ?C�Wc�$��~d �� ::�>��q��!Amp֡;����.�_���ۇ�s�R���z^�6H�۾��CB �._R�&��AJ��D?�/>k� ���4�5������W$����_�����՚�R�_��s�2��wX/�'N��q�c�=דFؚ�wI硎��!��hM�)����8��=dv��.L�)X����Le�][-�r>}�=}=�Ϳ.A*�O�U���̚:F�X�'��y�/ϭμ��y�O�8t*]���,S i;����
�R�S�X��3�S�,@�D��Q#�GT�-\\�Wm⣧��f��N�6ϵ��	�F�5+q

PI�z ��U�?��F���1 ��ǲ������a����)]E�g�R�n������ '�{qy���t��z<�:],.<���������u,|r=D=�/&����_�krjMdh���l,E�R�W�o%ny.���0��N��1n������F��"�y�G3�Md��w���b7�ή_�~����%_w�����/ ��*+	�&������Kۢڴ��Y� 5�����$@󧴩�s�v�:@�5���]�	9�GG�,%5*�р
��C���\*�<����1�Q��W�y	?���k�w�Wm�)I���8d.SyN�)fb=zP��t��NNO�#⟌��<m|��6��4��>�K�SݍW{�C+9�41�������Z���L�>����2�Gg3���mU�[�4���;��F�����b7�p������k��0�a�[|�l�zkăM(Xl�' �#	���;C,�#�uuH�S��@���*���`� �Z��~O�a�b�^h����ϑ)�yw������kuw��N%�Q�W"���u0Y۔!����8#�D�%�=	tڊ����iEŏ��k�䭭��< 6kf�
�G���'Hܟ 	�$ǝ�g9�9�ޣҁ��ܚ�b&�^aqk�5��f�X��Dc���_u���x%*����Q5��;�g����&D�$<l������fƊݻ����-.��&E_W�L]D#�C��Jc�~I6ß����
�ۍ���u%�V ���]7�gbǱ B��!�+�*x���G�ڻn�7����n|z��/p�{��1% &�嚚U�Ö�Is�i8�ӈڛ�J�wޡ�B�V�fƚJn96̧R��y�^)[������G;^R�ՌG�'
��6N�����׵pi��{���]Y��8����*Kψ�H�6�k+aq�7�`
R(�}�슧�i
a1l�lm�����Z�[�P��l��\�"\��Qć��6�:~��b�V�d��iv{���zb_�4�i� '�xFQi�-3F�bZ�i�h��.�HTV�"VQx�԰gp�12�(c�n)���`ٗ�����`ԡ�lb#?:4}+�N�`���c.�ՙ�nr�y��x>?4�����?��.ϱ?��UO�'k��v�����ݱICÅ�����<��t�p�_o�`�3�z�u�S�
<�_J)��}�d�~�Ie�Z��G�y�H�;)���5y�Ɋ�n�qvG@ȕ�q���{����O`H~�uX�xQ�J���]׎!T{M�=4b1����Pӷ���]	W>�_5J�U�^�۶5�cKj	iZF_�M�k&u�M��-��x�B	��X�77��[�z�'sDF���#�dG�d�&��b���9���l�wA��i�F���:ه��'���B�!�J7����g�Ij#ڑ<I�~W�g=���O2���?�ſ��<}ӫ_�m�U�*ic7�����v9�=��a�{)�t��?�1�u�{�>�ULt�p��꒯D)�Q^]0A�1Q ���2ǫ-Kṅ��!�eI�t���.,���`~����{�r�̸�x�$�<[!ʸ>�W71&NZc�ݜHCC'��P�ܜ���N���UeqF:=�])��]�°Bw_�D�����GW����7�*"�5#�������xc٫ٕ��s������w�4���g{i��A޷쎣,��'F��t���������E����l���d���Ŵ���R���R��7B$��o!��K�r_��B��hX��y�N�/�t�&���d3% �'] ���jڽ����u�l�=@Y��湂��h��PI�������(Q�<�����s)�wx�Dz�Ĭϋ���6�!�寣pu͋K���$�I����6..��I:|==c��,wX2
3���Z!�T14��&�>�~#ͷ��7��z���<��ض��P����� ����Rk����s�迈:c�ڢU+�N[�͇S����O7����h�pt�U�D�_�3��3 !Y��s�(�~3[���������[��=,a�{$:0���3{�v{v?�h�0�dJ"*�WZ����=�k
J�}��"V�_�I����b��2����焄艄6���a��a1L��B~�����:��Hߍ G%�{=MM-Y#�"YE�7��f��l����4��bip�/"�q���?'��v��x�T(����ܑ �J�u��K����}|k�9�N-k��{ �ը˻�����
�G���Tm���.Q77���� z��`r��;
!Hs7�5=���3���YX���w>Nȋ(�dI� \����M7;�R)�m��}�fJ�a>��;=?$��=
|ܕP���ā���
"Dm�wQ�"���h�޸O����(�&D�eNȘ[@O���x��M��W!�|��)�m������D��$����GH�XY��E�/�Ȧ[`/��V7�w;�Ү�t�O�.�gcIlk-�>�]�������27l��Hw�V[d�e-*�]�ؚ�O��~hR�v�!��Fc�$�Uԅ���ŕӉ�����SJ�]�7ozG���9xw�k6�|�n�"u$XU|�_����O��DFf�8�$l�-s�$5>P:�.���2�ļ\�$1�K?���Y��a-���N`J%sNA�M��q~���-�]�'`���v p	�C�U\ �(���5��1Sv��Y�i�͈D�{!�����e宥�U ��2�ċ��a�JcJ��)�L{,b\Z߉���ǯoV��T�s1-J�ޭ��/f�Uo��o�)�P����;j�0\�l6X<-�>�X��Y���HV�����)s����P�G6���0A g��7��ټ���03�iW���6<�^���fO��g���Q`��eT����|�d}��.@���ڐ.4Y=�*	)���I��Ha��=�Q�Ġ~�`W/��a4l)�Y�}B��ԔE�~�����_��Ԧ��e����Ѡ���3>�|��^ʴ���=�DF?D��W����3S��lE ���Pڢ�5��,�t�^I�>^~���G�u������ng=T��6n�����y��闫�(�EsN��ns������y�Q��� ��xl�T�8��i���x۞��*o��@�7����jXxX�ڑ�����W� �B7za���ң\��2��G��8Γ}�G���E����"'�D��Kؓ1ruu�ٵ讚�vw�.�R�b�6u�q��|�=�un���+���		PuZ/�ء$�.�1J����"�EB�W���f3k��̽3����gC��K@+EX��.�bx�)N_����'��yh�Ac���J�{l|�负&�mMW��#�N�Yi�:OJ���ք>�vC��W���\h}��N��Q)���*�U��Vf
mѱӼ��N�u,v���*�K�<"��*
Q�N	#E��t��'�A�Yvl��h�	Mեwe0��uK*0�v֢m6�uZ�����{i��YZS���W����g����VT�6�����r[
�RKQ[�B��=!���7�Ԕ9�N"�eD�*��\5-��I6�@$��\o~��;�##�4��?�~��cSa��)?��,ྜ���fZ�!ȝ���z�9��=ɿn�kwռO�7A�Cб%���~��Z��^�2��{p�[g�hr��I�|������er}�q.�I�w��~٭r#���ECz���ju��x��x�fj�eh����!9�փ�xy���J��ymBH�1&7��r��< /&�#��x 4t^c߮7;Y�\��Q�rb�����~�R�,{S�A7�%󣖗5я$S�3G�m�P�vf�o]y-��3��I���~L��Q}	{]��g&T��t�*)�?w^��Q�qW�%%R�/� ayZ�!L*?��G����o��&���S�?B�>������:�0hZ8�1�,�lw��=�<�f��oH�ؒ����1���hư�z'^=�r��Suj�sr��*\@����:!��dD�Rxހ�}��/<vf`�44����~�A��wo�Vv�	X��K�Ʈ�~9����E��}� �~�΂����e峣#�	N2w�V�~�u�)͵!9�*�7&�~*� ��d���"��*�^|�܉�]<�]��x_S�����P'��)�/���Dk�bkQ��C��:d�.���[�ֻ�����z�-H"��h�&�q����qD/�/��%?l��2՗��c���O����嘐f�	�n��T�Ks�a|�0A�l�K��$�M�=&���"�,�g���͋zb��><���۽��:^׳��w�+����)��n\�x�\����+g�;�EDF_�|��y��=���h�D\�a�o�X��ٶ�o���r��Uv�R ��)�CBZ������K�)vs�j�=�"�̈}w���q��I`؄�+�!RtΝ��|	%�T�*�70g���R���OXM�T�c�$���JRKPS���a~Q��!��g��蓦�p�c�5�xW�[ғ0De\�.��d䉈q�	��՗�dQ��G�k4����}���^d�a��]Za�>:�o�ul�5]=`����C����\�l;�:���3����8k���.����q��:k/L��1H�ߞs�7�ډ���N7��C�=����v�7.R� �-�hZ�z�#���a�`��2���,�r YO��x����4϶���y��4,��Y�Ü����N��\�_�2�6m/y�{R�z|�у�F[�f9sg}6w�
m��m ���	zů>cͭ�;��R��3k���`%
E���
*K!b��
��7�i�.Fg�G�=э*W��3z}�f�dC��Ko)*�	��ӻ̄�as��* ^2(�b��Zx�9�|�B�9U���������o���7�`�����'�5~���[�w�b�9���}�xp̾����/�$6!:N�N-�e��|y�&�3����W�c ����mx�P}���M=�O�����%��+���0��M������~�:A��l��gDa}��F�������o�����nO��c�"7�n����l)��/W)>w�Y��;k��
�G�O��4����S$~)K4�]�-Z��a�)]Ҽ��Wg���0��h�Ƀ+����04���Ę�M�����y7ET9Fݧl|y���bAH��;���Q�����Я�:Ȃ!�31���
���'��M��#�������6u��.8W?p�O;��Z����<0���.��TMx|!y��;:�@ %+�8!v����NӦ��<��7��w�D�7z����B�,Ao�4k[��2�s<2r�m+^- �!��w�ݑ=��p�Rq�g��NwK�����YY��|������`Q9����������-{Ұ����ӶC��:(���Q<
�zz�,-�=���6��u��-�B�{�P���[%.3>��㺑W�ϻ��Th��Q<����j�H{�
[����L�2��P�� ����h�ٛ��[���(��z��Q�����yJ��7�`Lg��m����͊|��O�~�ɟ��9���L�&���/�.�?��L��[����++��f�G�"Í?@�'"���6E�?��1ߥ�o�鐧����7��Z�f��"���F��QZ���|Ml6��ɲo1f��Z_��gV�}7A���0��Z�c���0�4vY���@M&0gԜ*D&��B����S|!j�M�8h�Ӝ�=��:I�kI�`zU�PM�mpT~T�-��A���E�Y]�)gC��V��/��5lь��I�_d�{��;;��ws�~fK���蜷��
��o���g��L��p`��wH����	��0�ż��Y�6ǯ� N�v�<2;��뉊s�	��\�w���0�vK�o>�k>��!�ӎ_��+C��}��S� �h��F
5ۣ�Q�8��m_( ��(�#c(���jY�H�^�� ̓����X�$@D;X��W�g�\cZ*�f��8h�������yB	���d��4�!Llũ�?e@	�����ޱ�/�$剞�,�и�4�����QyXi&A��c�K�A��� q0�OU�Y'^Ql7�~��Ǯ#<��b��:�������]js)w���`����I�@���n��3�}�9�n0�Ğ��N(��UL���(tp+bJK�Շg튈��P�יG���4�)�9]ʞ`p��^��}��:�u�_��W��E}Y3�X	h7X��r� �NU�v��aƱV��}$����R�B ���g������t}��P��P(s}�}�>`�s�6����v�\ʁ�y�2)�\� ����t�&���ι�<)&���]���������/;��~�Q��ϝv��%�h��AYU^�,O;�Y�\@4C��IC��q�ƢN���$V&�zG^���F�1=�D���5�ٴ/^�PT�m;|�7�}�P���e�0"�XQe��!V��|a�b*�xi��~��]���6׳�`�/����qؤC�"����	�n�}s��#+w{f��AT�z̝.EE^���&���A`L@����,C+�Բ�<�B�������m9�����;YQ���s��-*�������+�(���M�n�aW�?�dzI[$q� n>�m;��w���w���V�ԓ�q�B ���^�]�88�W��Q�@�Ϸy��Q��k?����^�_�h0屃�N�}�˛$$���[xOO�X��6���v��yf�y�����,���(��s��a�����>�S�J7���z3�ߞ'�/X;-b�J�;�u��G�.��:�W]�l�d2�_ނIP�;c߂~8�ʐ{�s����by���>W�hr��j_n+ː�.^i����W�j�n�D��L�(`���2&�j��cW�Q'ٹ$w	 ��q���&Ei0f������sE�~l�w��3����s0�6P0�{��#���R?��M-b�1�D��<�8�C��M`��A�Sq�8����"#��9�N�ϰ�@M3��ޱ����w�4�=ג�LQ��n�T��'�̊),���d�kj�dx(Ά����>k�m�^
w�5+�.v����C.�~N���������-i2{�ངA�4�
-�p}�x��G�����7����x~�񭎝k�%棝Dg�p�W\��Bleܕ쨗�ad>�T��*��GC����9W�QW/��W0��I��cDC;|�~r��bt���%5�h�.k�.�3��;��l�yPC�{>3�G�Y�d��~��7���3I�����Ƙ�T���������s�Acr�)>��TVY��s����)�-R��;��>%��8L�k�pP��31�,�,����	םJo��(p`�g~��'�w�����F���g�^�|x.�SXb���ޫ���}��Z��sb�%o*q]ڻ?�S`��+:�.	���br�bG��'d��$nL�E����[*�U\gԬY��ˡ�WpN�"���)��U���5p����b<;����tZĸ4�N�M�����Waj�W=u���f%ERl���-��MsZJ�gr_���&��gd���]Φk��� HRPV^�yl����@�����Z��o;;�G���͕�=E�(��LR�M�|��亝�)��5�e��db��.1���� c]rc����P.	`����BH�T[�����y* R�`�#�
Χ�t�Y|�z�I1�ag��#��'Ɛ��j�����#S:o�Ui������*�w�/�}���#�s>#����fv��5`�0�h�n4���=7J(^g��_y�	�cX~i(�Iۊ=<����Ø�6��m"�t����;I����B�UO`˟.��.�����B��/�c�������uբh���D�_l�>�P�e��w�]#:=���voF}�S�Y荺�ӣ�� @�!�u]��\����U����M�����j)B	 �%%iL8=�*��#�������ZV�h؉Z�FZgᗿ�4�H�Cq��=��A�PlcH�PO�?ѝ�	@W��o=��a�^�A�	۳=�fGҝ���>k��c��J�lV�bٗ���� p���8f�V��߇��z��	5����{�11k|4�UBx��[>��^^wFn�Du#��UB�qT��
�'�����}Qx0����G���J��ľ�	�k��Ȯ}��'(��\�`k�������#(�:Ĵ���v�2���V��	�(�y�϶\���c]/������%.n$����z=��bOk����)�I��$���)��X�f槎�#<4��~'���{[}�F5������z-R�ד@[��5l��:R�	uz�Y'�(1����Y��pIXKC�yFO�@R��܈������^���.�����|_�:,	���-��>T�j�,��<W/���޽��p:�ҽj�2}g����g�V-a����8Y�)���Vp�q�Q�b�W[���3b�cI{���k(!��,Œ+��߃�����*������u���
=���!��� H�1�P�F�l��L�$&���p|�b�Զ������[�6[�A�.�:�w� �/z���Uߊ�2��������V<	9�P�dK�%}�O�"��A�`ۢZ�v1kKKf�����ObA�|DČ#�\��y�o�FjQ���������O�\�$����T�v�mz�D�����jC�����cb%�s|�_.!kR�����ʨ%.�F�3�'B�5.[$��bw�/ϳ�I.�����mKg f�,f�����Fç,�4�
;���Y۠� �A]���J����N����%�N�����{�2�L��vT���
��aV��=S1S���Kؓ(��e?�Mޠ��˶���' Ċ>IL��R!�R����$ҵ(I]XVQQ�С�n��r~������z��o鋢�V���J�x�xr��o���2"�&�?}�����(���h�8�Xj���4,�3͡�.�<�:��x_Id��I�v�**FI��w�=�Բ�q�����T���GHR�M���A4�cV�>O�e-��	�FV�dX��t�I�(&Ϙ�'=Z��:8�`��_�fRo�K���.����yx��q�����qi�{�K=����,��0��޺�͋�v�Ҧ��aE�٬����֦�Wؠ5���_	:�B�����"7n�U���Ts�Mc`�?�Ċł���?��N����fd�	���x��-$6�Od���z������[���������I�B8��n��`�w,����S�dr�M������5Fm^������64cX���ӎW/-��M����Y��]�eR��2��C,�\���z�r�^��ddgT\��ʯ�}J�b��~)�0 ��'��Q�&�q�q�޾���4��q����ǌ#|CV��/���nW��r
�G�w�{~��������H]�.�x�v��Z;�E.�UT�=��ϼ2�H�0!P �
��̓X�ǀ��ÀM���	��w	8����v��u<�*|���zS���9�<��a|���
S6�w.F�{��w�z44�C�%a�+ũD�1�O�I�h���������7d����e4��%�u�}�_2RR`�z{�����L3zrrr�a�b�~E�������#H��m��F�	ԋs(�9	��X�#e����r�?�'Q�;��'?%�m�bI�^64J�Iè�B
k���VV�z��������÷.)����� J$�?6�*���w�x�<���)�� �n����3Ͽ�ȏH7/�t�����>k��.@zŋ�]�)�������P/Ǯ����wa��]��cIM�|�����nםw�j��)Fx!���Q�tk˖ �!Ȗ6��8Vl,���)�Jl�j���$��ۓ�83��b�@-C��H�8?~��x�K\�X��K� ���	�q����nb_�,�6YZ���Skk����!AcT��2�K�h~���1�]���oj���]"�E����ra��ԧCW>� ������>�.�{`�!;�$�{��UY���:�%j���_�妙Z��1��B���܂��'����=�Kq|L#���(��}���S���6;�Ӣ�P%��ѫ�a����F<Q�0`/�:��#i�r\��F3S�g{��O؇#��_�X�=>*�2��MX�B��P6�_��O�٩��z����H�r!������*fkl,c�h��Ty�|���F��j�jz�׾���L�2Oͣ���SQ69S!r����4ZZ?��>@��Te���fi)��m2a��z��ýC�W\l��N��ן����Ч)[ b�����zT�--�@م.��\
pFb\4�*��z���E&��e7�[�@9m"i�.}���a��%N��v�3}z�N�r���Et��~���`��~�*��7�����Q<Q>Y�:i�S3|2�? �,/
q�����j�����t*	��������v��dW���w����W��u�}z2�	#�{bcD�q�z�9��-%��)Wj<�+8�j�֢��^����!ަp�X���.�a�x�G�*�Ӌ�~�Ć�a����<��fG�8tRUXt�$�-�"4���g+�-]>���XY�����:ZF�Ku�K�u�����SG��^�.��J�Eẁ���'�2�j��][N1���?���Yۺ�����*��j���B6�m�\.����OJe��w���)a7�uY�8!3�こ�P��#��_���On�)x���-����޿���ż�hk%^�����e7ld�N�$~3ɪo����:�$%�y�T5?$1��ؿ�*�ǈ%<�Q�&��/���l)_�Zn�Lu���E�2���J¤k�����$�'_ߌ�e#���w��-'�F8�i�N���w9>��K�ƹ%��eO���)�v��yv>5V�$]�(��,�̤�pz��¢5"67-�H�*��aW��o� B���kG���+�7o]�ik=��n�>icvM���/y?�L��cH�,��&�M`[�I�1�� u��G���@
��5���by����Ū��L&�ys��i��'�qzrN��.ѣD'�EQ�e��C'�Q?���5��Ѝo���g�t���㘃���k��};j(p��&�[O/�*���|7��<�e�=w��|�r�}ȯa�L?ć�Nh�����淶~pt�A�ߦp\��k�؆ʀKP΀ː��}[���t1�C(X�\�u�YG[;y"~�ts�Z��K}r֡�U�6�O����[v��$��ۓu��b�u�����9:����U��_j�~�-"E�M>e�%V��*��^�]���*�<�U�Z5�H���Ю.�R���w���c�W�c�������x�>_��G�l��dN�� Fu�
�=��@m�?���V��)�2�2�v���3�Ye��I�a�'QW����p�
��*Z��$���K��-~vk@R�ISH_X�C�Ne l�e�S��\�~��B.��������Iڏ�T�]�~/A�`\FH҉ۭ�>��QD4�/8�o�z(���f������e+�;5'�ml!q�5m[�L�=Z/�C����OՖ�UL��s�x<J$O�3���,��?S40��O6;�Li�s�YP(����9�N^�(��@��U���V��L|�s���:0� ��ux���ei�Z_)�7J��?n�q�&��ZVY95f@sSTb�^����\d~@��u�����M��Qg�t�쟻���t+Fv��e�%vu�2��c����t���D[��BI�J� ��x�XM�C6��Z;'ViL�����t��~�qS_�0"��1�����Ϻ9���j�1�vĳ�,�t�����t�,p	�9�ߔ�m�=��=�<�N�ߤ�>&S��0wv"#W	c'�]��tښf��F��UW�ɐ����ل��@@A�^DM�o�	����z�^�66�(V�+�̙������}h�k9�/6�6��gh	wfk�ŷ��q8v�v��ቐ������P�H��G��
��Ȭ,�������^P������O��`/T�Je��`Ɖ�q����N�ǣ������a-�*��АTչ��Y�Ng�ўV8��q�-���0�ʹ6�LP	����]TTF5Y�rt����]$[ �H�rDgn�P��4���A}<�*>�|�6�W��z�G�k7����C���*v�>[{/�+�[ibl��K#$��_��A\���}�O��I'��xPIcg��0��UMh)�!�qC~,�^z������b����m-|��o�
W�8<|ChZ��S���Kk����FL���<�Z�V�(��8e������,�7UM�B�5.k��H�'bag�T�*������$q��#�i�5�+��
�˥�M}���R@K������m��¸��0�lw�BI)RSk�~����z�&Ѹj̛���&Ufyyyy%l<��D}j�n}���g��L|n�R�!Ig����m]i_[��޸���[vn���_��%y��䜜?dz]�r�J�Aq_Ų%3p�����/.�v�����F��8-w�t��(�VU�ghM�r�}�38��:�7GK���]L��x��KS�4���
�����ze�z�'��z#�k@���=��M~<����蔹͓��W�k��%-`�O�؉϶i�K�x�Ƙj�����<�._7�!�S���H�ѣ���h|Z�s��<��_�7�>x�����W5--_��i�������R�E��w�Oo�L���e�[}��^왉�:���w�Ag��흜�I0�����,��4��<�u2ܾ��S�ı)z�LW2ļ��hν�m��w��0���,�aKz�Yf-��Y�,�b� %N�P���8�񘍁����z��*��B"<��ò��y�US�1X�����7��0,(��a�$ä���6#�1�ݶ��V>��
�z@�uL7��C�ȍ$���I�6Z�G*�"M�y��w�2=��ʵ�|�{�ħ��H�P�J�"�#���6�1V�\�r��^:0B?�H?�37������+��ݯ|�[��^	�L����������A�Oǒ
������j|off�ں:bh����_�7"s<\\��;��)�l�Q"��X.BE]\���8�13;�g��;;�gdd��&6FN��q�|����^����A2�T.��Yg[f1!&���}�Ķ�r~�����Mp���J�C)pGe|����q"`&A}�9�p�qd�,#�Z�MP�0ARa��e,' ��X#�"��k�얦��v��QJ�u�����v�@\�ʳ���-o�fQ	��21�%b�v>EJ?0)6�~*��2ݸ�X�x�F����f뫬�?$�UX[]��E��www)�R�݋��[pw/���w-�w�����<��E��s�w̽�"ۍ�&N%�0h�����*+�Ư"I)c%���9�"t3�!��İrn��Y�d��r`M5:�hg͞�jm-�]޷^�Rt��b�k^;��Q�bPXQ��qqN��^��3�LJ�ѡ{BL�Bkq@������l,��t����ʗl2T�Q��2�g6VBÓ��»ٿ����f��[Y�u��'G��unSe��Bx�|��f���,�f/s\s9[����ׯq=�3�f=�e���}���A[K�t��H:Q���jèBS����H�;�� -C$!^���]�ԯ�9�����o��DQ�L�8�N�W�=A��<t8�R�^�i����R��1ֈ�TfY�O�}�o��:{	/�^����z�rҊ�u(�#�|e����j9j/��Z��&���p�B����ph��&AW�/���9S�8'�"��[h�/�d��]�8��Mbv�m
G`����C��E.-]�!�Ɓ�}��-w�Eoy;mm���,�am���z�����?X\�\^��6�S��K�gxLs;<h��5B��ѫU�5�>���1��,qxX��HE�$T��H�(\��q���V�C�N5�����ɟ�[�����C�y���˧�Čhc>��'R����RH_4	�Dj��pEV�1�C��rnbׇZת��|�����[V1����5$��
�M4GX��Pf¢QpxP�<?��w�Ye�)��aC���ך��<}޵���l���*����T2��u�8��9K]1�d>8�$ƿ�oM/��`���I k����U1�`�R@�p��b�,�ā٨yNV𫒗�6��rIT2�I<��h�:_n S�Zz��8��eɴ^y���CV�қ��I;���*���1�V�w���Ѧcn��r��LXR�ߗ"�d�{y�d�oB�%�\�J���ȡ&l��UR��4�_$	�9eM��g�^f�9�>���t{�u�2v:P?F��oxo�W�Y��>��"n\�p�k&
,���ÛWl�����+�&a��T�43�ګ�7WL�H�H1�h��)p���Z�ܒ��˧�O��n�R��u���T�~W�C��?�����О������UHf�Jw���k��Bg/�s�P6�f�q-�۫p�<Qk�6+?Z��<�b���m���Btmxyx��r����
�����g��+[�,(�*I�!���i�"<sV-���\�X��	����e���`���Gr�Zq>%��C��%��Q䮥˪���_a�����6�r�;T�����6XN7>=�j^�ɹ��x\����[Z*���T�G}x5k���*(H{��Ls�=@��J��puZ$z���b�qJfEzy��:���h�Rv��!N�@��� [�ӂ��$tR���җ��|�-}
a�Ҏ@�[�k�Z���t6景��*�ٚ◦x?��D��8=x@�I]�7�|�sx�W��'�$���{5�=�ٯ�`U�(���4��n��.�LV�Y�Wʦ��[e����A1@��f(�f?��4` ����&�Q�$�fq#���*)�Y׽��0���"��JAE1�G!��QeI2�b���e�4�N��3�����(��~��U��t57���|�1"V����>��[A�}�^��������_��r%��se�"���U>l���_��fD.G֊9���Ύ�s�����~	\ԧ7��ѥ��:d
�]�@\���gu�˥��sN����l��%�rMH�&\��2��It
0�!�O�~�
�Ҿ�����((<N���n��W��B�7+�={�O1q���쥯]L�=���n�I�,�.���2rx��(L�r� �������+���HE�"���Z�uO��h��$h����z�v�9����P^X�ѥ߀��4wK��q;�����������rmg����=�#C}{]��K�S$	.#��ٺ�}�cP2����=I�ꪎ�~�
�[Z�F8R��m�q���+�����������t$ ��Ͳ�^W��i�B8{G���`��@u�tH������B�"���\	0�8��c�рD]Nw����smjrU��:H�3�cQ�<����Ze������Üev� ������.��k	��$
�d
,��2���b�G� i�a�����l?��<|�!�*(V3�r�y�lr��p�	ӎ�'���f��{k��Y=Ӆ���:�㫳�=�{�WY	b�����z:����&tlJR(����^Av�s�(�ѽz'��6\\���B�ʡ:����cWِd�t�����.7��Utd�}�G+Ȅ�Q)�ױ�a��bb��jj�ۣ&caY��k{z<�bw!Ǧ����3���CCp�>G��.ii�4ѴC`={ ��� BM�O�X %��o���[�t�d�M��ڢ8{ �WRh���.d���%��z���?�L��22�"��/j	�}������5��Ŭ�(�R��b�s�����WO\
����έ%�E���-ץTS�Vw�1�a�i��#�R�/rY��Xw�A\|0}������q����"i�R]�-2�/']��Y�z_EI�L�^�di��>\��Ex'Ǽ�E*��暈OA�H�,�MV�*��'z��3���=��K�<�8ꊃ2�4<��+� �d��ʆΨ��LM:ƇA9�
�"@a"��|�u�i����!*<������l�9����Ѕƕ<�w�=�t*X[^]���Z�L!i�
<�H"O��<�>^��������x�i��P��H��S6Y���f�9��u>�L4��p��O��H\WrH�=2��n^K!�Q�Kl�;p�*ᬻ��a��⛀�(d�B�Z�#M&�~i����L��1$��fidN��D�E�8D�߉g�S+�������8[g��Jק�9J'�J�z�|�g;�s�D��
��ϡQ҅��m!`AA�r�E�&��8��A�(�-����r(4��}>��jna������-s���\B����2oP�|�^�+��h&�\=|
D��011�ֶJg�H��%]=Y\�R�XÚ�͹_~"��Q��b՞��2�n�������g� $qn6�D��\x�V&���<�~���t����&�3�]�#D�*y��.���x�]��A��K�ó���x
�
��4��� �z@�Ccm��|��~C��^6�~���3��
�����<���|�2&+Jݢ
&��<�mj�.-�3p�u��"����3��;��wӺ��q�
�VዠY� ��O�-�����	�¨�F�_�.O]91Q&Q)�]��t�}f\����H�����'��@)�E��!oZ��j�B�.m�S�D���?���(�BJzq)���Q>�Ŭ�V8��\��,_�I�#�Y`�8����#J���@/�k��%2�S�)�ݦ��H~������I��	OB�ؤ-Y�_r8�wK���g�:̨l��}�g�ڃ�����/��)�c8f��%��f|�Yq��J��� ��&���%-��MB��fh�>�Z��>Kt��xߵP���zu{�:�l'��7&u����H?(��P 2L�� q�Cq�=
A"�6QVx-Y���u�a	8�v��5[�20P�xGe%?�&�i}�>7{�����D�u��C�mo�`,-]�\��׷_�ZmV�@σ[o��?��:���?IQ���������v
ifڇY��P���Ê��;�h���@��xTɬ
�M繶-H9<� O��Uވ��U�"QN�d�Iz�KD�ç[�d?����p������w�6C�H����o��!bh�2�c�M� �����݊��J��H�ξ�M����	V]���旒볥��k��5��I5�WoP?���xȲ�d��D����Q��|i�ip���L/��B[A-�v.5�g�&��m�2�Ӕ*�0���eE\�*�����������^H���B���Ę��d�;���Vԏ
�5��8�)��
ʘ�Ÿ0A�
w6��6ω��yQzUu�����j4�X;����>���"����zR�u���� �H
7GL�/*�B�݇��Ӯ.��$W�(rR�:�,������F��1 ��:��Xt`�����o�������~g�/�ġ�*�s�g�8�������J���"8�����N-���E�q��2.��+M
m��џ��>��a���e*�ث-LT��El�u����/��zB�3eΊ�TBW�%�~$��&*t��3����rW#�8��ͯ�)o~��h_����/|�U�!��#"�X�2?�� �B���Q,����d��(׌y ,
�,�jk�J�%~��,���NN ��3փ����"LJ�f������C�x�!!�A��?!���>.䆩�f��7a@�L!���D��\�1ZNI�nF��L�ǵ\���O�̤4��jq�|2%�dV�3v�H���|ɶ�`w�d�/�����Tz�^Yq�7�3���]�n�#O;M]p�٤�X�I���
̩�oµ���A�W��P֘��Vi\��W��c�P�	#���tE/�[�rc�I���-�On��kO�9�G{��
�z��t�w��'%�V�K���4��`���#�%%Б+��E8�lqC�����4�*��qT6���*�?��7�"h�Ĕ'�7�p��3�-!M�o��B���͆�f�#.A=��,r�!=�?����Z�o��[�(A?�d芟6s���Ww�n�!���,�q��
4����P���<�'���@Y��^h�r�t,	dx��=��b_[�����c��Cd\�8���IJ�T�%�D��IJT~	թ묗ϱ<Mi�t, ;<�4�&B����U�l0%</ k��-A9�ߝ������4�~0���3ıKS:%J�R�r�~țG���!�
@s������9�>1(�)�q�K[�"�X��u-6��!��ѵ
�Ѫ�_�<;�j�]P�	D=�[��z�5�mj���#�x��qD���l/p,Ev�c�yE�wa#c%#�m����	���,����ߡ�A=Z��,���jҦ�|{i l�µ�`1$��ݹ�l������I03ƈ�|pH�J|׭�י)����k�O
<���Gۗ�2V(���@�n�E�d$�Č�pHf��γ*%�N%�.,Ki��mL�o��v�͞s}]X-����:��Z��q�;8B�E�&�!B���2m�T
2[��v}j��I-�q�	��X��vpJ�����T,C�������M����Yd3�>��H�]넅�C�����M�C�,Z�s�}_y$I�klAn�G�4.�"@z?A���M���O�78�`\)�B��Ɯ�z8��Cd�Rp�WP��Y��qh$zb|�Q�4�
��OY?iϣ��;�)7 �|��5=����n��,xxtx��"���t��>�+}�j]�Ɩܭ0|�rG>�� ��i����J��u�f���?�]���\VwL�)���C(�Om8����g8�_��[���ė����}��黩��{� N�cL*H�w��O��r��)S�������`�,��.���P]��jX��~ҎǁV�h�I�H�7�y|E��vE��oc��3��9\#O�3�C{2��3Z�'4r�˓�S�5 �묶�ljP�xU�[q�#]���uE������˒i����mhJ!�/8̄:��؞�y�~��$��C;�R�6nǖ_֖���!�M����.�<���z�z���obZY*�ęB��֊�0&k�\񌖜Ե�����w=�v��*�
��|�9��A�,�3ԠO5zYՋo�ɯ��a$�J#9�EE�_ ec��!�x��%�G��S��N����ʝ�g*We];5���0U27��s�~#WH��z�kBh�q�W�^}mk�[ڨ��)TТ���.4���q]c���<$��Iՠw���{��qw}�FFψ��ˇOA �ƹ�2��S�@ ���8s�m���'S�Ōb7�-�7��')x*����F^��I�+j��E�Ά�m�!�fQ��;�ٚ�)�4�e�6ٔ��&��tG�S�.�ڙSȣoȧ�O�np;����H�?�c��C���Nm�B������?A���N� ��'��S$�ƌZ��)�8�S���׳�M�4c���SXH����w�cH�2��ɽ�.�v6"�Jz�%��"$"��{O׆��a �t?=��՞u���w�3�s�8d܆!?4�����mn�j��p��	��QI8�V������o��3I��<�x��w��Y� aG1e���g
�pFe%�̜;����z��w��.�v8QByA�3�cOW]�t!qdj�vj$+���m���Sr�1$R�6��g~�oG^=����n��2�~�r{'�������e�3�Xm��F��%��D����/'���l��2��UNr󱚌��]��f73~�����7l���$m�)�Ú�6)�g=��	OxM�Y�s1�:�7��x1���x��o}���u���mv[oo�^Ef��ݾҮ]�����t�J)�6��2��xЂ#�CC.qL�E[�)ݙ���[�`��d&�x̼��h�*�C��BI@�WĄ�C��2Y-�����@���|w���6^����{CqӞw�ljw7g8��76$	.�+��hz0B��(G�^<�]��d�Ӭ4��g�<n�[��j�����wjS}��x�{�̴����|};#R�D"�TM=��
�X�nF�_�[9��}��:#c%-h�*z������-��L��ga?C!2Kg���ã�^�����)�[����O�f<6S:�*!Z���|����|�?
��/���Pf{Pb�  b�E���wi@��Daؑ���a�T+���4P�X-�Tf��&89�U%81=::h+�0f�a���$ђ�v�l#6������R��$Q��	z���#�`*�WU�g��D�;L�M�t��(�$f7r�(�s�""Gؘ}����t���8��mUWj�W�١E{�ޘ�^����])>�	�7��?�J��-fCf�Os���t��m4�IK���sZ�I}h��i��ꀕ�5>��������3�BR��k��2C�����33<��9R$�NY�����Q����9�L�O:5�,	sKC*y�7�o�t?YM����d��%�����)W���N�Z��AyF8�0���������B��[a���y�>�`6�v�h���6szd*R�YG߃]�9���ˢ��.�~��Y������䞟]`[���0%n���xD���1����&]5�Y�؈�p���t�K$�V�rC��Κ�I�Sl�[�F�����G}��M���t�,��e��t�/j8��Jc(X%^r����A�2��އJj����U`=`����s�=�s��T'bmK��~����2��&�I9 ��Ի����Gz'q�(Uu��ZO���<�1�Wq��j�p����᱿��C�����g)x��� �ÌH��vt2>n�4�D�=>�������J���Q��j�������Ų�!^:��g�
d���
Ck���Z6��0v�����$�s�sMƦ2���R�ջ䒘ߴ�k���nBUi"��B;Ga:C\�����	m0(��Ի p���4l�MK�:)��������)�9�i%A�Yeeh�CA!�<X�Y�h+��v�N�����z�𫯒�2ぐ��m2u��̏&�����|Zm�!���	~j\Ü ˯}��*�{�d9�k��LU<��7��1�(c�\A����B��:GS!5��4�,��g������t�[�v���\!#x7U�T��[W����{=�=ܾ���R��zBo6̬}����R�ܯ2��<��G�b#@���-&N�8���-1���N߿�ḎN���R.#ꅤ��+i���ވ�նN�?8Y�ӕ�K�r:%%�	���ͯ����dj��|��im�cQ-T�6quE7?���TM�I�A������T�$�H �=Yq���Jȗa�h� ��l�O�k�ez�=��j��`�@�Z�j8�Ь��M�җ۝�~V|��+��7�R���~%���@"��Y���5��>jô�ܜ<���=ىμ�!A��D��@� D�B���V�ƠV$� 8��3���i���14��yZ~<��F���ޠ;t`�WbO��蓝�%6�R'k�d��i*�̀g����������W�Hm�ÖWL[��P=�����Ox�;���`E��̰ד��?��}����&�-\*�9�/Ӷ�@0A?��p&��wqpQ!�&2G�#�+C�����e�m�US�o��z�����j���؟�gA�%������(�"ĳ��� ���*i��o�.����_���t��Tx�W~g��afXDc�g} ���ըk00iv�LE�Կ��~.$!��6��N�{A}��3¤�w/�7e;�2�>6*T����u������=�Y��E� lu��;�9F�@���^�ހ�]c�3���l�$k|��(U�Tȓ�٧��ݎؐ��J�1c���qG��0#Ֆ�_2�,���1m��^�S\=����*�����f��$t���)�g$*���m�J������;&���}ΌyHN��v��\Ԥ���¸����q��4YH���"�:k��ʷ+h�{Z4z]�:`4�WBNVz���ē\U��Ii�n���:���&�c�R ���#����9����h2{����ds:m�=W[t��>�{JE6���N�X'���p��ʎ��P�d�B��X��k�N%�;�+��MH���Եs����ŭ}�n����Ҕ��4_�i�i��{v�*���om4[�n��� "��R��y����Kn�wY��\䭽�l��Cn��z8�Ǹl�w�͞w+�iEe?�}y�W�;
�6׉��&$UV�z�ҥ3�u�(����}�|�>��Mج��lLa�iD�Y�e6�K2&�6�,��qEI@�朥&*GF�������-M��S3� ��!>y7��|�����|"p�߷�}�I��r΁����� �Ipz壒tf�;���jl}33�ط��<��7U��*c�I$?QDʇB�inD�/~�>�({�U��Y�K$I�|��v[���^w��ɻ���9K��4Kb�Ub˷uH�d�P��G�.%����Z��(Y!D��ae��@�=f���=��HY�m�]���ˢ�0���HC�d1�ˮ}�K�{��K��R!�Z��`
���k��u���c�^�^T����R�W4,�>��x�T��?�oV�!�%F*3���50'3'*����y����E����E��'T��.bZL2��\�W��qlf��n�c_B�d�1�����p|#��W���_���? ��ŕ�Q]I ��j	EkVg���}��N�W�!v)�&%#𞖣�r�m�x� ������Ǔ�^����
�Z�s���/����k�8�d���5y�2v(#�����ܮT�$A�(�򟝊�j�˷oJ7D����A����ۻE�SN�"[6u U[8�HGۄhh:K����"g,I�8�l�A�{�����a��Y��U����88z��S����/:_�wo����Qd�"�����ll:��@�ze�X�Px�8�>8	���b=�i��~���3%_�H�a�U���K|N�~k��n	����JQܬ\)����S"�5?Q�b�#�v0�
�0-��. t���3:-���SɆ7����?�4�m��?b�c�Hӆ+#������?������&�s��͕�zM�^cY%�2+��Zm��5'΍��75!��th>�L�tl!�|�}���������/+*n:냑�i���d�Β�M}������m���tCSӠ����ѫ_�l��ڟ�lcvG�"�� �&mP��F;��=<���Ȼ���]j|U$�9qg��&;v��ퟠǜ�A��_q]��+�b1�(ܴ�8�1�KQ6�`d������r�z�����ϝ��c|k�E|
�W[/K��o�^9@C��/>���/�&L2^({Ia<ϛA.�<tI��Ѳ��OI��k�1�4�/z}V��{�'�LH�	9�oo��i'NVb~LmGP�fR�XN%@�l#ƴ�D��+�*C��.��k歚p@�ܦj���LT���)�$P��S�k�a�xV<���v0YJ,3G�%p�����jѡ&!ci��2h^m�.ݱA�0���xȚ�_і�ə����YQ��
�Ӱ+*��n)"��U��� 9�/O�vz�0J�����A��}'�شX�̆�?Z6��5k��q��=jMa/h��`��|��ٵղ�Ģ"E�삻�_���8`*c�
5F�X���Z�2*UII8d�L����!�z>��{k)��9,� qV�d7��8ʿ���i;Q�M�߳���Çd�С�a�i2�Yf�Q��E��c��*�l��{��5�)��:����<�Y{0情�	��'�Ľ�xq�Sq�QmdL�w�3xR�?E&���W��X|�A&���Ȗ��X��M��oN�B�J18�s-]���6n��]���Y'�����RM���c�Y$�?�J���aY��}�軳FZr�lHY��8�`�=O�hj����
&�[S�����8�bҏ�MLM�\�����|��o���`$�����̛@��z���UK�vx��X��ُ�^�盃//���ޠ��;6�;�r�ޕ=��56�|tcݾ��B$ZY<{�x�E��w 
C�����$�xI��n�
��g�-\급��N�G?�#)o$]�����GY e���S*�sij^�������q��U��
����V��E�Ȣ�#��
Eh��A�� (U�������ԧJ�M����*���P��P�%�Xg��!S�Fhz6��u��1��r�N�D^�>�=~�f��LG:�o�������E�ORt0�����>�-<.�>���*��������J����=��K�����G�J�6�ͽ��MJ��u�5�{"�M�݉n�7���쩻��!�<���>��cS�&o%��|ENS��y�����9|���e�����7X�����0Isq�h��R{��9K�R�Y�ӿjXrI�A�;jr~��v����KC���B�������s��������+S�Ew�7g�������ޓ�E)bU�����g����Yr��O�$���$%$@�l�hh��j]���V�ֆ^O4Z��86��n���yO�~���6 �d^��F$	�3RY>
��9��)>�/'	*�)�t���Yw=l�:���gE��1}��zb~x�X-U�l��ߵD�yr(�������ݝ�ֽ��9h�	�a(Q����5�5�^�x*����";��Ph���~D8RJ�F���}������o�jd�Q��ʑ���N���7��F)!$	�b�I��ؕ��ڝ�H�S�TSVY}�B��(�cݤ�C8�>P���Ņ#�
_$f��D3W������[j�bD�C*X���x&u�H�g���&;.̷��;̻�$�f��B�Wz|(ҳYm���:���;L��Z��8�+y�>������x����B\��h4�`�uձe΁GJVU�H)M5������]��7�\0@p6A���ܳ�"Z盡�Tl�{/Ծ�%��E����d���!51����H��ԯ
ь��ŵ���T��}C���p�� (�ٺ�mF)�U_�+�R5�s�7�\�yn�( ��:�ZqeLf}kj`�|���������*����w+A�c���[��������⼗i#4�pb͊��>'���Qc:n�hZ����Z�-���:v�w�1�Mn݂ ,'u��, ��ﱩ\������Uћ�E_�Z{�5��J�E7jd�����"�4J8�Η]�ֱ����2�9�rAB��摶�8���u�aoV�[����t>$����#G��$y�������[�D��u�bx�:hj'a#���4�
�eÝ�~��۹�����������Y����g&��y;w\5�X �oSQܛ�O�5`�1�eI��U���s�V��㮚�]��IO9FU�Ȃ�紕�?�����؝�]�$K�����S ���«:ْ�"O��F+�8�i���rL<���׭\�U�q��0�Qm��3
65��.?u�	��ƺ�0��"�f�~my�x�z����o�P䑞0��g( ���	I���hn�͂J���%Qn:鷷4ؼQ#����r0/��$���V�#��_N7|x^��='$ꕃ�,\7r�;�0����{�O�����&�`�+`)q�.w.�%���K1�����Q�_<l��L��&Q@��̄g��.��i��G�����'zZ��|�gS�h����>#������xǫ����ͬ2��n���P
�p�m��v�H+;���>�@`�E�hq|w>�߁��7��%�Ԧ&�XV<�����&$l�-�+Z�<!�ds�t&K;;�b���yv\����1���
x���(����oV%)�Ц?ߢe|�_*�Ƞ^��5!��xi��7s�[����ݮ%hؗ���!Fj�z�"5p��S�Zq�`�	�L�*V�0�(A#�j6��j�ѵ��ū���I.����2�A��,������$i�XuZt�+�\��.xy�a6x��-�-���V$��fZ�R�N��3�b�|/ H=����7N��6u(ĕ�yT�>�*��
�9!�#��}�v�@L��k&��܆^Dbc�w/H��QD`*Hzn��Q����,�Dd��$}��%���]��CE��r:�x��z��xw�����T~G�U��^�g�Җ/F���3J����{�ӻ\�Us�Z��� ѲM���W�p<��0����Ӛ]�Ӵ���iKC}��(j��LK������G�'�5���>U%A�� �,6���iU��@Q +)LJ�A�^l"Ǹ���l�b�
j��,�LY�ؿ�W�����������'����&�^��cִ!�8�XI)
���y��C��9^���v%Z�TM��i��2)}�˽W/U��h�Ա��>�rB̾,bjYW�{v���{�Uy�U�>��.aڣ��G�LS\�}5�*��K��I��I0�vl�S�L}�2a���&&'��n�jz�v�-V&�R ���65�-�����R�<�)����_�y��s]�*�`ջ���;��D����X�G��n
�D�A��λ���EP�cP����Iob��-�����`q_�qϴ����ƖZ�i�f����u
IQ?��-�Q������c�%+�;�$��������@!��Y2=]�l����糞x��;V��`���4,�:���:t���vmczjي�;����L�[�(�Ե��-.~���誹�]�-ݑ��L�:�����9̶��.2K�Ucb���ZB<!D�}�S��R��Wq_��d�ɲ���8d�� a���P�����]�4X�K�Ā�ఞ��؝Ԓ1��ޢ�I��2[m:E��V^icvO�8�p2��D�e&��@�+'�R��g�b� 2�-mc��+Ma��x,�jPo�xD�^-qD8+>R�Y$��Y�S���8%�����v�����5G.�9u�O�Ǻ�TK���BmڿT,���na��8�債%7�w�r�WYс6�dL��}��	�}a���mԑ��Q1W`rl�e����
�\��4��2��~��d͕;lZYibo����������M�<5��c��V
v��{��,�N�eP�O�XFC�z�;G�oⰫ�j���V���š#�KǬ(�&�t�M�*]�
���3
����e�$c�`G֢ddZ,�����{t���'�%&����}��5�b_:�	��r�i��Igd�abe�k�+�%��(��L΄ͭN���4P���)r��F�!��dc�9ʢ�#��;5�#�Ԛ|��}�R����[_�"���������PdY��a����w��Կ��S�˯�ҔN��3?�h����I4}�F�%#�cT�`�W9��$Mq�u������78�!8w����/H�u�A��^��6�7\܇P���>̆�c��yIe ��)T0�o�7�f�İ�� ��MUu�!��d���[���u�������	N�e�b��Aj������Tn�w�\ ��;;���Č-��c��j����T��.��<�wܤEre�������F�����nv��D��+�Ȱ��(^ts�eb��W��'Y�%l��W�^k��Ώ�8i��n�Cn�H[�D�����7�2�03懷���f��j���}j�!輶��c���CE3�0��m��{"�Pd��ԕ*��Z����zŃ�6�C�����U5�/�vV�n9KD��gf�͕?Кf5s*a1��]S�≩'>�� ���M�M���'��'(����f&
� r"���$k�r��*V�u�S���W��1I��3t�;�m�p��;'F��)-��nW9%�IemJ��!�X
iI���3W��,n�٦Ŧèe��|۳���������Ql�-G����k߽쭿7��P��W�$�HS����q_���>��{����k�x���т����.��{CWW�=���}�
�I���)�#��\;���r����c�b��;��kz@�\��0K둙`VR�ߓ'���ʖ�J���`O����>?=Jϥ|�I��k����u���H-�sO�)��4�k��+��&����t�����~@�
cDR�Ӝ�����P��x�.:5e�
-Tr��g�'?��"|���x<�x<˰j�����ӯ���y^iU���FϪC�I�Jt���깡���⋠�8�$�t(Z��|�3V�6>0��rx�~�d��� i�^��!���a�>���6�C�0����y�ш�=��<ЗA�,�Ȥ_����sd��n�:�:�#�NM O�ޔ�w�n�W��}?g��F|��ba��d�y�K���W��t*�f��-]:���n��D��"�f���ġ�M�O��iv�{��[�9�9���n'�x���l];�j�w���v��[��$��Z��R�ݝ�����2��!/�H8Ɏ3Ʊ�����]]~ז����_�_�Q��X�I �_̒(D��\�_,�ED�)�aw���lC�U��oDE�K�~g����spGԁ0j:����ztD��v��#!�����Q-�����C�^*.���x�&��'Q> ����E�i��l3T2dƈ*Pc*��LN�5���AD ��ۥ�#�Kq�����R|y���%L⥧����6
hx��@?.�$��?���㷡-#�tW�Rk;G����H÷k���.�,@~�J�Åivm���%�_����n�����%��GW��&�9�\����y��}�/�T%�k�p:�:��X�1ߟm>\N��n��?TrI���mr�����*ML}b�<�e�(�O}�l�<I����f������)�/3f[?���Y��c�j��c%��b����J=p�����z�i��0t�7|�3���]����O:�|�~I�����OҍH�_p���5)m��qX=��:��!�,q/��xl�P������2��Z5��E��'+��㧧P���w[��������5`v�L��5�\�q=W:8��{��T��I�fa@`�w`�dKJc����+�d呈i.��$oQe�Br�=�� ���%
��.cM_�k5N�ɼِ�S|�C�
� ��H���w+�����*a*&*E����#�I�i�r��"���+#/��K��k�g/3{��p��/6SGt���c�}�nzA!��L�O#R+]��͝�I%J��L��i��h�N�Nc8��%?�oQ�}O9��2���5ssMp|LHr�U'�2�VI%���ٶ��lq����1*Ymm^Y�\2YI�:�vx�\��V�4��a��?f����(E��y��<A
k��7�]j�<��j���i\@e�-�XClw��,]��\�K먩����ha�8	\d����*U����0��_�����ѐ��{BAY'����!w=4��;��'g]?I�c�d�W�1$�ߖl_�N'�XǍK;D͢���ȓ�I�%$|��Ҫ�����pǓX��e��J%ZKMGŇ�^���NU��� Z�}����yk��<(�d��bG\ےT�,�)Qd�I�.J�6[����KKx�%��)���d.��	K����K�N�L`0�똱ᱮxm�\�4���q�e�V��p��*��P���^;)�E߽�l	r�M"T���2��4��[�6�Y>�I�nxj�P7�b�� ��]i���.��Ҳ��:��A��NƉ�8�����ų
Ϋq�u�����yF���b�����=Vddl�+�sZ�x�>���n��Q�5��+�D��� {@��ɤ0O^�'����\K��@u�n-�����5!*�R���Kk�9z�nVv��+_�S��gƎ�.w����/�[��1)��<w��!����u�yQ�$)��!����3�#ՒDJR"��ѩ��:W�y��hj"������m�Η�Dڊ�N�9r�i����<q\ ʊW����v�)���)~:PD�|DU���|^+uoJ4��$B #���\H��&+:I�O`{���ՋT���c���!=k'^g���'�� <Y����X�jv��C�L�~�]Y����?�^�����ax��l��e��V��}�C��n�ha�N�Ga
���.O!H�!3	�I0�Nj���<[kq>�PHe�� �& �G�`kk�k׮q��E._����&UY�����277������tgfh��7	n���4�� fggY^^FOF�7X�ш��mV/���z��pH�$x�F�ʂ�;� ���Ci��v�!��"MR�$�3�c���^UY����Gp1"���^(�m�Ⱥ]~佼��s<���\�������sgy���B�%G�8�ܞF%P�궩��*s�֜{�5ξ�*� ґ��L�� 0� ���}�Լ��V���� �'�F/�C�s�+�vhP�E�rT<�[��6��)~�1-�S����_��\E�6��>�E�\��.�����y��7�nj�ݧQ�T�4l�#.����m�87;f�HZe�曯ҿz�'�0�hE�Q	BЬ��c�{/������s���?��p�s�0���^�*sbQ�4��/|�ؿo?�s� i�&:(
-4
���$��-�$�H��8���p�H
����#BN��6 k&z$�h�Q
[Ulmn2���z�
W/_A	I�3C����αcy���%��z++˴�-H��4�xL��#x���U���(�9�,��&�9���H-PF��TupJ�#�D�zd������)����1`�BKEt���������U�
���>���!�y���>Gx��GY�R^���ؾv���6�;vr�"��)NJ|;c�����=^���ZG;FDY]�x��Fc��j���
A"�(�Q���D���*�/hei���1i����T[��Ȳ��Lw�S����ЧxۑJ!�j�����?�<:�4UN�5��@���'1dx�ԙ�.l�Ԑ8��
d�h2T�C�p��.~�i�.. �"R
/���j�y�Ï��曬��
���9���eǑ��{�A.�ֹ�q��?|��n=F���ؽ����������Բ�¢$�(�dH�Q�Ę�l����)$�R���Y�i�ı:��!�:����p8���?�W�Z�t���0��\�em��5E���()�	�s$��چ��We��$M�F7/TBIRm��޴��������r2�6��H��+K?��ˊ�=�,,���?ex�
�=�.�}�]�|�9ο�*	`҄�~���v
&�0h�
�c�l'4����$k/��m��lA&�%0T�=���&u��.��Tj��P!"}DFP�
�]-E�d��O��^�|�"����������}�����<"���S��ۜ��x�fUA�"�z�l�z�X�p��a'�ջg�(�#w�%,ʹ�=�hD�(����^��������u��\��`T:����#���9G���L�~���Ӑ��+W8���� �罏}�{��n6�C�Rĉ�N
��4�4��j�n4�L��
Eͬ�=�VfR`��=�M��)J�	��C�,J�w�}w��>�e�`0`8R�.]���1����'9�n�{S6g�b��*��!eQ�j4ie��HO�\���E�h4b8���j�n�0J'�QMv�"Fb��j=��%{R!�����8' 2Mx��qN��&�ٿ����%^|�i�^��c�8|��8e�&�ۈ���¥�������>�\�J�� 6�[pu1���a�2K�c�sv.��<n�C�L(SC��:0�%1�-I��Ea����ޥ+�ee!/�U�k��~��m��/L;�)�V4�`T��E������Wv��^#�s"T�&<O:'B��Z�(E�_V�L RC��v|�	%��ND���X���s��wގғ�_
��\	�ՒC�y7����O}���,�ū<����o0'5��ۜ8�J���ݏ����E>�˿ċo�N5�*kIS�H'�r��Y��H	18puf:���yO����;DТ�hO�U��DKI��-�!��s��F�/�f�,M)&��F�!��(��L��,k'7!��%U�e�M�bd��q�#�mE�� �@�5Y����
D ���'N�#�&1�X;�Eo	.� >֗��W�����Y=��f����
�g���/]&�)3�K<����[��G�!=RH��d)3i���op���W:��X�ȥ�Zh�B5���6��J����!/��1��F��v?�!
"'��U�
��R���$�n�+((z}�����a���ӂ>�ۆ��}��<��D�(�s�m��,�\���1$EY;�!�A�\ H��J\Ybc ���iE(s�0B�����0��β b���S��q+�މ-�(�[��h��W��?�>�.]&?��V���x�ť%�~�c<��WХ��|�3�/�_�,w��~��5����0��NoRmh�	��DkISM�ۢ�z���8'Ѫv�u��Rib���"� 1-F�VT�BjY���ZvC��e�=EQ ��,�#<`�%��zb %�V�f�IbUU1��U1��� 0YzS�fn��m�L�p>���~B֗�=HR0�q�cCm[V���k�t�ۿ��;8��\9�D��������w0��Z9G4��HR����s��˴JG�� �	݌�]{i�'okb��j�S�J��٦��	�a8 ���u����('2-5�Y���dj
c�U�h@�Ώ#����_�Mn�G��q��9ô�O����D�H�(p�a�[:��enɲ�?���(�:�<��`E@��R�c4�h���(�p�GS
5o.ʚOW{���,�Ho�"���f��~t���)V�x�R�,�?��y�7��? �,M���?d߁[x��{��SOb���^`#V|��~�~�C\Y�����K����R�b@h�8�!K���i5S��J
�VTUI>.�*W��I���`��?���ڤ� ���^��c�yd�/���Uus��GHY�4���EKy��^%E�'�[KU�x�PJ ��P���b�Ru�IW3�C����B�%ڪ��)���'D�EU���:��Kt�[w���}l�^��_f��E3kr��G�����ܸD&�4M	I (�Q1*y���?<�r���'�?�ұ�d�w�!-=_aff�E� J�3)U��.�3�|��B1�%�Х��zp��DKP2�CG��U��6�����T�1�6<�+���쟿��n��/Lw�S�-�3o+�$z�D�۴�C{gf�N���� "m�Rxʐf�,Ck�N4i3���Z�NfQH��h'�NB�u�^J���������K/0~�T���U�qxd�$b����~/w<����v����g��u¡ێ��dia��O���wq�!�����O<A�iS8��U��/�wG�I�i52滳,��3?ӡe���*�J$����I�"K��}EIQ��G9ei�>)��M}w�e4��>��v�,ͨʒ�`@>cmEUU�yN������ں�s^�9UQ+��L�IF+Ii%i]�儘�}�u�h�R�(mEQ����ል�M������V#G��g�����?�vT�e�ʞ�|���Hcv�qQ����Z�!� H�J4민Ƌ�5v�v9r�]�����G��sVz.� ����X+�F�����C���)�5ʥY��Y��]t�&���0R�-$YbH��D�9����']���>S>��_�̙)�}��<�}��8.�S��)˒�P����G5j����\Wy#bS)d���a�6IB�hb��DR���*KS�('kk�X!�t �v9q}��瞇�+`"^ZB1͔h=J5��ct{�w}�S��^��o���@X�������{� {�G��L�r꥗���!�Μ��|�w>� Q+���*����s5�OII��baa���9�mZ����"�0�f�he)�,!5)j��0�iu��&F-�M�Z�c�F��.<�2����UQ�*��,EQ0��F?�-�������H�(i*C��b�ա���&AKu�@'�2����Z<������~0���?���Dv.-�wa��,9����=D���ˇ>�I��u7�҄$A��-*8���'O�����N�p�#q��'�� W���~L�j��-cc��k*�������J�-V�69��ŕ"g;�\���6tn݇ܳ��!ˀ�5#^�l&�FBKK1���������Q�\�~����_�)��)~�0�O�GCք�"ϑ!��*�7������d�%����-�N�4Z��8(�pH>�	^�]$l�����>��b�$S	"z��I� A���$�D`9mr���\��w�񩏑�H�-e�֑�%��9��>�)���zcv4�����ڷ�{?��z��/1�S���wx����������>���뗮0��$�JD��� ���h���lf̴;��BUZD�����
��d�s.��P'bM$�a[U���6)�d����x<���~#��F�	lԻ󲤂��O3��;�f��hM�&hcj��jb�Z���Zy!J�J�UM��&�cmX�A#k���Ȯ�p��.�r��ER�!u�]w���x��:l�Fac��l�
��m��/~�W����~��﹇���]ɚ����A�����[b�]�1ӝ#���g�_��7��v��HW �a��a��-\��p��>��@&��,&s�,�ͪ�a��y���8�(E�����)~.0�Ч��b������R[{���'ZYco�Za�d!A
U�l �sbY`L��U�UYa�����zOp<�U�:�k2^�YRu�>!b	G\A�9���l=�囧h���a�E7��^�M���±Ga+�)#v5fx���g��K|�C��sqQY�����u~���o����tM2�"�f4*)l��;�`<f4�m�т��&{�������^^���ȤD:�r�LJR�Qb�cm�UQR�e^P�sʢ`42�>`KG�ק,�:�H�.���41#Y��L3Dز$Q�n+��i�Tb�@�Zy`�����Z*�b�ecMt���B����ê��i���|8$�%��&{gf�񞰱���st�AD��;���?F�0K%*I�A }@'�ܗ�����!�=�>��O�������Wxsc���F��)���l/q��x�{e�νt;]�����{��Cs�;$���tf($���$����)� %�y���]m����i=�$�9"<��?"���z��1������/3�}��()kW�ʂ]�ܧƣ��{�J۾ ���WHcj�Wሹ%�y�G��L�4k�W��K����4d1�␡ j)���Gb�8R<��h�{<����o�!��+��&�[ra	��Z'U�W3������#��_'d	qc�[�懿�G|���}{�!��V���c\<~�?�'���q��m�]�C��`t/�X���('�O���I�P���I�S��f8�c���s���MiJС"Vc�F"�#�N�2�h�2)��IT��`K��I�6j��8����DJ��HK*fӔ�$��HL�H��#��2օzd��R(b`9�JG,%A9��c��W�H4�f��N��Dr��rD��p���_e�k���w/��_c�[Y��ap�eM[ht#��7x��g�����Ҏ�����7Z��x�@ـ�=��,��Ǳ�e嶻�3K4J0Z��̱���<��ϲ8�WI�ÜF��=��%� (��S:�i���;�JF>�ϖ�g����|�eESN?r���a:r��'���"FF��!�=,�/�h�.6��"ACU9BȤB+��X��"K1Y�r��G ��3�'�%BD��]���ϓ����%5�@#v(ɵ���?�<��%���Œ��Dj���nk!G���'ȇ�<�����	�}���[�}��8-�qY	��Ͽ�2۫WXٵ�d��v.�^"؊�Ը�"P2�VG�l�ʔX$D�F�l��B��h\2�6�C�U�Q��4�9	C��v�P��	����v�C@Y��"�z�m���C��� Cmx���Q��(�ѓ�.���P��a�k�R���$al+���(��T��=���������ֶ���I�ԬW�cw����[�����B&��N���0�A����5^�ַ�o^��t�|����Y��j�� �عk��b�@!X$���2��q^"0��u���eL��Hf��3CPCP��^"���sM�q�R�=m8��r��\x*H���������p���/Z�r��Ę�)~bX0�&EU�Ìs����L�T*[�eR*�� �h�+R@tU��豶��_�@�R
�u-�
uX��?z �-�U���Y�h<��W�Jsy��?D�A	|��*GA�
ې��K�fh,����lT�lty�����r�}R�h�>���D���y�Ut����2�]�׮����i�n�������s4�&Z@��#�2d�-����~��l�������1�ܤ�k�DM�qe �BH*[�R�DӜX�FW��E�aU[_�����u�X�PW�E�	H
�pB�����ђ  �$�կ'!���N�ݞc%�a���W�ظxd��՘������0�6\0tL &����v���np�$��~��;v�|�a6�\�E�4�Q9$Q�V��*�QJ�C�+!DM �DL�F�*ٱgǿ�T}y)*��$NղH�G�����m!ŕ��D>�Ex%*����,�ϲ�� N�s���g��6��$"�D�(t�G���Gwg�,u�!8�4�Ѝ��Z\8p�Υ�l�xbaj��3�5{2��4�9�Bi�����M�E�0��ŉ��}���$J��9epM	��?����Z��}�c���� �b�̸��3���_A[7��+<��{y�[H���ϑom@�6'j���2�w�c�5O�E�W������P��b��cR���ع8��b��vJ���2��)*�%�
)��,S42IjI�L���4�e� M@�z=�%��eI3y�>�*PU��*)m��,��x�^ �� �^E
�-��b
ϼ4�nv94����]T�9��>��lmW�����`���{���o`J�"�%����sM������/������ؽk�+׮�]�ck�'01�IRD�D���dT�(�C� ���ckK�Vfݫi��"ӌ V����^X�R���HL3!�*����֨����	A��E�p�3���	����}�;N�#h����U]������\�gNJ[��*MfB8RJݴڄ��ԇ�Qz�{�\�N���&o��E� $$�0ڦeRv%��U.�ɟ�ٵ���c�}N�dD"I!`�.[��������d��p�_�)n4d~���ǹ�}���O���d{��=������]��p���6�p`e���st�-z�g��%���c�F�eD�	--0MCj$E�(*A�"EUbm풗&���-|�%����cM�df��DIS�4���!�}=M���y��("�{*
&nsR)B�-�r¨`!�8�����y�&Vva�/���h dʑ������un}�{)����i��a��DH;H+�����6�=v��عL�0Ko<�t�$JA�,0Zb�1;yO�l����b����Ο=��kK��d��3�E��D� B��%BF��֑)%6G��>�x�C/c��J�F��:�S�aZЧ��c>1���nF��u_i�Z	i�ۊ4Ӹ�xL�&�,�,J�N@���^�5��D��7�K��qj��bHBA�BG�"��r��<�Μ�ܗ����Es�HYB&��B�[ETl!�����יI�<��������K�������bnn��K,����~/�9�k�gi--�gXy.]�B���-�]C�. �~ںz�`���yE(�[%A�z|�%!M��#����$�UB	�H�c'"b@ƀR�>�(�BN���9�C�`/-�-ɭ�m� ��s���-�%4*�H)(m��Y60�lshi���v���a.kp�C\�x�Vڠ����᣿����n�V)$��]5BKT�17�����m^��r4���	Z`]I�m�[lth��Z�u�"��v -bPS'�#Ry���6�b�3Y�3Ϡ���鯯��� �ރ��D�z�n{c2Q���*gO��]t�ǚ�/y�N�*/1&��g?Á�.}�#�}�+N�#��m��V�w�1|&��P[!��Pz�6U�H�V��qN��Tm4�4�C��6Hc����8ѽ	!�����>�]h���W�D"uD�@&y�y�����d����1�w8�hT��q�Dk	Z���:�����Myu��f[:.<��{����۹��1��滔~��� �%K+#��׸:ڢ�Ϙ�i�iwh��D?/��$^ �A�G��u�>TDFHd�	ƐI���~������O�6�!L�>�F�����\��X��}�eiUEn+�x���>�Ph��<֗+b���UE�s2���5ӡ=��&��!W/��s�Y��6����d���`4���,i�fZPU �@	E�K_�~�/���e�bҤ��[�f�R��q���	v$ۛ�\����=��~D�1Xw��h����x_r�қl_]E�!I����ĔYB%
F!���m�@�jA����K������?��8)�|U_������?�;����dN��iA��Ǌc�RT��T8�P��#�*m�P2
��iȄ�����Bj��Y��#[)��mL�od�#y�u�JC$_��]�i.��X��& ��n��T)":TȪ"!eA6�![O>�r��s�F�E�!"hҘBT(+�8|#ᮏ?�O%��_~����YN4R���^f�;�ނ�س�@'K�tu���7�_�Fsy��}��G\���z^�mi7�t�M�IB��1
���e��J��s�o��'B�S%�:��OϴN�QPY���]�琄)*G��͑{i]�T��_=��y�����u���EH�j�L�Y�����7�֮r��5�"���Ҝ[��'>�;?�I��e��s�3(!� 	�|U����_�?������}���(��Q]�J��b&m�ѳok_y�1&�(����_aa�A�� d��N����O����5��:\�x��,%I4�p��E2�(IE����*�Y����+�03��i���*inT��f���b=�X�EI�$sf�<ŏ�w�?6�y�#H"ò�;/�w;�� A�o	/|,k���ĉ�5�f��T�Y�1�Aw4gg밑$!i���%%EY�di�uOPG���D�7;�:�4Ȉ���F@�@��T%Ki��~�)��f��A/́�ز@�a�(IQ�����8Fj���ƕ7�dGw��Ù7Oqj�I�����i�;�9����-����%v��Awn�~�G����`#�i%)��.�A*�Th��!��2B#kzv�<L�W#u�8�n<x1a"�j"3��Ι�������9��y*�jݺT�D�X�����b Q�,1hi��=����p��CdFs}�
�ш�5!MH����~���?��i������(��V���ƒ("i#p�k_���0wq��Z�`����4���\;�ʾ�eΜ).T8��iF*1T��}�������Tk\U���"؂�_b�aH��r}���e�c�	Z�y�����t���IZ����!fRT(��Qn �}�P*��ч˾r���f��y�{��՟����ӂ>ŏ��,>��ۇ�>� T+3o9�0���d��i�9���F� �#�@��N�sH)R��B�u�}���9O��9b�_�.JQL������#�C��,5�,	ɩ?�E�����!w�Bj>�
�Rp`L�`T ����OО]���q�ě�Z3�Z������|��ev�����<3�׹��f{{Ȱ��8|���,���{}��qemA���Y�f��D�V�Ƥ{��	^�;n!	R�V�12v�sR���ps̞Q��^6ĺ�ԗ!&�o��ɔFGA+Mi%����n�oq����F�9{��k���"�y;��g����!���<'Նf�RSO��ىŹ�������c�J��fQ�1A��UJ��5�~�Yn��'	yIҐ��"D��!Q�L��#��4	[}��m�rǠ�bNFt��^bp�"s����Ӗ�fWnb�E��,��	�H�Z��
�0��hfL־\��vh�A���2�,i���v�S�� ��d�)��8���,$	�|�0���Q>�����*�|�Sk���W($yUҞ�����w��#Jkiwg�J�R�z��5\
��6F*��	d��H!j��M�=i�A "AD����@"PAQ�JR�D�&�t }���n1���,?�q����4���;T���Ր4U��)<�x��_�_�������zŐ:{v3��DU:�q�X(���"��	����U�`4�������>�L3����k;1�&���5�<����<ϩlEj����ݹO�\G՗�H}Q�B�$Ww��$�i2�z��&&FB>&��m5��i�6	[�����3�*d��l�������'>�΃YJ4����d�&��*M� bIt%����?�C���m�U�Q�p��d�M���v.������I~x��f��2��0�ic2�H�bX�0BD�@"4.�I�$��V��M�ktƁN� �W,e3HRڝ9��&k�.�
9?K�]`�]A	�e����a�q�5�Y�����Ouj�/�������(��&{�t�G��/�iA��ǂ��>���ш`m*m�������;gwt�%��Yt��o�_��@D��eY���q!%�9��eQ���E���I�a��BN�7F�D����\M��ŹʡLF(��;.0K��b#5t�O<���(1k�6�U��H����9&$2���W�����/�L+D4�(����D5�������4Z�4�������Q�����Ć���&�~��,�*���(��; �BHA��¤	B��9�[UX�j��d�Q�����G�a�w.��P�ΙoR��*a&k�I�(�k4iE�"��Qo��vWBLR�I�q˭��c��0��b�g�*&d��2B&��K�s��_����Ӿ��^���]`�����o�� �fy�_�K.]������;>�N�~�<T�e�"�s�*�xTc�4MJ�*�Eۀ�,]�d��izg.�9�V�Ԟ�V3;��m�y�2�P��A��M2��Rg��ׯ1�Ռ���q�H�9�������3:��@���t;M�4��W��s;�_.Lg=S��q�C�#�\I I�9��s��Ŗ�D[��IRT`l�(Q)1JՌhjb�@!�4�9G����b]E �'V�RJ7v�����]���fq�0���-�d���;5��ޣe@v3|ѧmR���|�.�9�>��޻q�����i���(�*�rX�o=������ͧ�Ⅿ~��N3�-+h��bT�~�4�2Cg�
�{����f���lloa��-11�����
�º:in\�IvU5	Hq��k��j�&�=P��I=���K� (�1 �$ѵ�NE�U��!A�6)��s��hHE#�,({}�~[�� 4��s������>��wM|����Ȑb�"Pє)�9���`�;O��?�]��=��� ٨*�+sz�!�<�!�ށ?s���?���uμ���`��zU�۞!��۔��y����XD�H\`��g��yv/,s��[=��Ƙ,�4��SbM���<FJ��Ue�þ`��{iwv`��C־�g��u���r����$�y5�DG�?��U㪤�M?����c�.��/�c(|I"��
������z8�:A�Jl^��#1	_��c���h!Dp�⽫=��5#] `�BŚ�&'���쭅�:��DD�dޮ�B�U@�����9u���c+�`F�_~�+J������E�����P��#L��d�(A�^np��>Mg�a^��9��ӌ/���f)��1r��N��y��f���9�t:�j6YݼN��V-�s�"D|�E�Jg"`���/�ʣ�	�y��_F$�ࡌ�'
h��$��PM���HP_T��l�i��$t�-g�h�	2xR��!�^�r��&&_Ib�q�����=ʞc��iF)<�y�W�B��NB ���*�gߤw����%��-�m|������w}�1���^ �2��/}��.`+O'w���S�O,�ݵ���=���T$Y�5�Q���J���ŵ��-o�s��6bu��mǬIh'>���b�C+�XHV�d��w�罏������K����N��ܤW4�)I�d���\i��1��H~]��V\���왒��`:r��/���|C`�1�Nh[ݽ����#{ˠ;����%���+��$J!�$��D*z��"�	1�ݣ�������i���|�Vi�����4H�ӑ�xdt��#�P��(E�**i���'S��f�١}��t?�8��KI�A�#ܨD
����@��X���l�=��_�S.��,�g�OK�&�lΖ���"jn���]� **�aA�<.1��E4l���CIl)hi���:^���`B�d�'a4�iTY��9a�F�'�t4I��E�=���f������PYʢ�	xFy��t�r��{x��c�}w��uq�ֿ�f�HF9d�� k7�%${�~���WN����F�Q�pT�j+��7�c�p�&?�ғ�~�Y��f$g��ͼϢ�D�SHK�s	�s��sm��XW��b{L���^�J�&���F�[2��֣�"J��2t�M2;����,�7P�P��<�-G������=��+4桛L�=��-��'���N��AI$�v�q�����d�i1�Ч��Pw��;�3Et�Iq�.�vX�ɕ$�H9,pѢ"���1ل�%�@&F(D��k%�R�Um/
��"�VY3ڕ�/��)a#Z�a%D��!#����tG9��_���k�O��w�\Y�G�"�jD�E!"� �
�$[Zf׎Ev�{��/��w���q�������iSK�F1d0�q�Ԑ��M��t�y��} �`󳳔23�5���TJ�rlAC�d���)I+U4���5i� �(WO?�DF4�QQ#�e������eM܋�&f~��ﺓ>�ｗli���F�J�GۊT%�".��4���r�������G]Yc�I����C4w����|�o�I��'�ﻟ�ᖏ/�sa�*V͉/�1ڕ�t��ӗ蝿��iA3�;���O'(VC��B�HtBQ�Ct��H��H_�T�
�~���*/�^��tY:x��ty7o��,��ۘ2��rc��l����>&��C�ym��h&ӏ�)��1}�L񟌍b���E����zQ|��lw�hLS
pT��(�"bB͜�1�ֲ,�=�oĠF���}#25Hb�׋��������ɤ]�:���]��
/��L��k��X]���� �:��,׏�����/�y�a�[:M*iA�Z��%Fhb�����%Y�îw��O��͵W^��w���W^b\���Jh7:h1RRn�6�	.kR9�M%��"�]Z���v/-��ڵ��S�D��<�@%!Ȉ�
LQЊ��6()Jt�������p��`�P9���XHMB��7Sf����;���������s��y ����7�A�ڂ7��I�ũS����W��Q*#?��c���ÇɎ�
Qs�Hx�������Sv���u� <�]=��w�����2�2��,"
��&�r��%FO�#i���)�0dH��$&�$1���neX#�"�J�L��ʫ/q��%�I��C{�}�����#��Ͽ��K��$teseck��m�|��%!D(����{���7~��u�����)���
�<*ƹ��G�Pw.*�[1�������B+M��7	M�7
q��n��nضʚ�'�*����+�QԆ2QL~���AL����2*�5�$<JO�G��h�M6��u���a�cf��a���2U�	5
�
�۔�����V:;�r�=�q���g����l�����U�����f�*��c��ۊ1�h<��-�$ ��j�#�f�Jg�`tJ�D�i73$�bk�j{��9@CTl
b������#�	Jh�ˊ��E�q��ev�u���!��e�`Ǟ*
�I�ke�
�[��4@�(!�(�(O��������ڟ���f��2s˭��+������Sn�X{�%.}�In����	�_?ɾ��ȫ>/}����ߡ;�q`~�l�'ɴB��V�:A�	�X��ǁVK�LR���1���7[,..����m�%��:����#$ж�w�*������gH�wp���t�mw|����d��$��v�Cp�ّ�Vd�>�d8[�K$i���N�?o��)������ly��Q�e��-d��f^�J+�u�HC����w�"1���ѝP�Y�:�Z-cM�b��.�7���^ĉ{Y���1��;"2��x����!"��R�"&/D���9-�^p�W9=�}�� qe	�5�R�*K��Kt�HD@�IH�fϞ]Ȼ�������ι~���K�>s�Kk4}`6wtU�Jҡ�F%�J3tE2.��8O�J�VX��2�2Ea �0p�b�	��Ѥ:�ɨ�X�
��@ޓS�����Xܳ�=w���w�Ck�KL��,���*�M:lHd�{�T�0�E
�o��}���_��K�Y���p��d����g��7���ȵAKf�ٸz�3O>��;o��&\�|�a�c�\���k�1-:
�| �b�
�QҔ��I)bI�+6�1���3�R UD�u��U�� ՞�t��H�V�i?���k�|�4+w��ʡe��F��q.��+H)�:T^��6�����$|+(�=�U��V�~����o����I1-�S�'A��,E�$!tC�R߱�%�`K� "1�7�nߩ�B�P���D'N�0Ӣ���V�����F�߾7+d"�F��D����Nֿ��CE�����|*a	�օ9��*c�jp��Y.l��W����ô�1?����l�h��Tg5�>
�. ����d�]��{��>B9���S�����ј����_%��u�ҡ���f�ei�&���
����*'�:��&~�Bi�L�0�����Ǹ���9|�I�fߞC=|��{h��ұ;h������%�+
�(*�J Sp1��C���|�:g�z��_�fm��s$�&��뾠�t m3�q��*�K�y���[��B5���7���{���ӏ��O<�'�`��W��il����T�$��&8ƀ�	�1hc :�8-)T$4��:��'R�
�f(����HSj�O>ͅ�_�<r�C��Ξ;��j��p��NR��a� A�62�0��x�+�a%�k�e��Y�&���)~N1-�S��F���c`�-��G}䊐�v@���Hc IB����+G�[IB�Go)*�I����� DĈ1��������v������!Pg��0�j_NQ
��j}��0�JR��@(�Qa�&27�*zW�ZAC���ی��_?����2��G0�@ʹ(dE���b��L'h�6�&Ah����V�-@w�����^Uǥn}�{|����X�r��#!'ll��i�i�A�3�1���q����(	e���.�"cD
���2w��L��5عw��u'��%���Pu�*d�R(�b�-�D�P�H0�4)"�T�l~�E~�o���E���O�[~ ?���/a��
�?�<�{�d��}��(�����v�*��.rh�N:F�����w�U��s���h6hi&)T���c�B�u�{U �@)���f���=;�<����h`�ftmc=-/�JEb�G�ب����=,���G� �Ǿ�[��+\�fE�y�R3���!�Y�+�>�_�A�>1|-����Ԇ3��C����p���˂iA���}�1d����P���������.�N��C�@�R���i.,P\�@g\��D�*CGH��1��O�4	1ܴr� G@����	7H���̿!o���MS!Ȅ�QKD��+�(1�AI��2�IA�	tJh��"�c��1�G,I�m���ml��8����x�}4�$��������&��;�����Yz ����rT�9v+Go��vxϯ�֞E����^{�8G﹏�#Gx���y�,-iXXY"�[�T#+�I��\3�Y}��s<�އ����#fgaff�����簞�j���#qB�#
č�DF�(	Q���M|����i���w���i:�.�=�({z��у�D�Dර�Y��ۿ��o=ɭ�x9�2�X�_�
�Os��?̑��^~�'������{�k���78���(=eH�llD≨��<��X Zj�P9� ��A���C��3��0,i�FI!I4��E����먍밚���7����?I��nn{�}l�v��K����2����h7����� �A�!�&E��G���>�9�S��ô�O�&�G�-*��?�s*� ]�IF)0	hC��$s�f�]���zh��!"��D�z�<1��%$_&�� ��u�Z��Bk��DL"CU;�����l���4
-�D_۠�J�yk�Z/�Q�=/�A�E��$�#i0��7O�u�2�_!;v;�}�к�.B���1qq�
���(*Uy�4�G���9Rh�NP���3�ڳ���W.Ѽ�.v?�q��n��i����q7�={	����=��D+E5S��Ob��X�B����m-y�ž�b��AJ[��={^�$�8-��w"
��'h���g(Og�ٗ�?Euq����}�f���Xb�+N�:M����}��<��?�4;�u�~��^ !����������=����i����	i��
\� E�B	C� A��?{��$�u������{�ԥ!��$@�$4%H6�f�9g��kv��5���1�O�F��3��ӂ�C��$�I� 	 4�
��RE������#2��6g�	�*K���۽|�o}j#�䫪G&5F��5�Xb�$��@�\�2h�h[�zRϱ��H��<�Ɵ}�����/�ݘ�ז1���~����'~����anM�,D��G��g��j"M�@)��w�޳�n{W˞�e;��O!(�F�&q1^����pn�`\Im���A�j��U5�Yߦ7!E����y�Z�p)Q��I[cT(�2�oݕ��$�: bPW���D�0-<W�|=��%�O�=w���K"��%��$T�%�*�ds�}V9�A�%	!҄+��Oj[�Ͻ������Ǭ>t?ûo��p:Z񈷸�G-�m��Ri�d�aA�N���0جmF6���l�	e0�_���׳��;�T��w5�ѿx��?~��~����ǭ_���e�	��\}�m;�ũc����k�2�������j�Q'�u ��)r1��ѦH$`���S�y�_Ξ#�������)N��*���e+�QS���4<��'��?�kn��V���QX�ꛎ��?�kN��In�� k�>�{��&/�ȋ����}�U��-��<vҐ�)"�_ZFc�R0hT�D��d"�m,�miCKH	kLFXĘ�*�FFtV�G�ºmh��w%�آ'�Q�|��0.����X���I���f�X���F�$���@i��Z�w\�'�ʅ������o~���?y�ީ�����-����SDU���i��v�	H�HA���-�n��E�0�){�����L���PO�D�LB�:�\���+�s�f�}w��{L��I-9���5���O}
N��֋�)d�A44�����L%+1s�'�D��!��u�m��!��v�zG$s�mA�gZ��#���4_�&�w�����Oq��؅���
�Fb�Yl�*�f̈́��?Gu�4�c��~�q�r�´p���Xz�M�;ŸF�:��EhQ�=`���4�I�vy��ѣl���)0�\s5Go�����ž;o��\�0Ih�/%E���M�ƀi,	m����J���9������X��be�fX��D�j�{���P�uE�][��gT��S\��K���o�z`�}��Il+���y��F���4W�5�o��â��"�kLf"TA��H"I��P�b	m i��>K���ҵaL��01)`�	q���F����	~� ��q�#cp�f^��w�ޏƲ��:�f=amX����\�����x듇J��(�m�����ZV��U��-�ޕ�go�.<�P%��F56�6�O�Ĭ,���nH�a�GcK�5�HL��PO�z�#1�b�o��6'EU:�vJ����ή�lISW�Υ���0.����~���G��f�B�s�x��j8\���8ߘu�!g ��	���y��j�3xD)R�	i#e�gI�N�A945\�z��kgx��O`�>��?Dy�}��}���:,�d�m��t�8�2f�5��6�����%����`V��vąұ�o���� ��5�ܷsםp�!�K�z���[[$��8z�-��яb��Y[Ҹb�z�7hah%�(�*րm�dLu�5��'��'���oR?������?���e2���
�����~@Zq�����[����,��xA���ޛ�����|���'���B�ʋ�����_�p��FC&q��)�3l���JK�N(�G� ���`����EU���M�./�$ 4][!�B���3��I
1��UE��84�}�	7�@�!��Øo@'C��>�Q��"�x�����%N`)"�[s��_�}1/���6��w���C\������߳w��9�={K�6F����b���ʽ�GhH&��YMU��p���0&���BP���uK�6c���*ٮ )��/��u�z���&�t?$�$�q]�!E��m�xq��(+��m��ZH5�����R����b��<Rfv�BW.Ȩ8������&'��R��W�!Bh��o����9N�>��/<�?����Y��V��v �/��h��*���}���S��h��_q�;?�H��C�P��+�a�J��*fa��1&6�P�_��T���/\�!�B��n��P.3~�#V(R�����=u��W^��8��	��J��͑�b�()U	�)='T����KKl�Xs���cl��;>�V�Ze|���y��O��=����n����mN��l����2�d�b
L7�,�����p��;?�bH��ɊR�g!J�<�''�N)H���ʠy�c�)�ڂ�z��$4l'���c`m9��_<ˡۯ����H�H�m&�-���QJ!�SV{�;�顡�#6�ӂ�ĔH�����/�g� �s�{�K���`!�L����'G��_E�ikL�ȳ�b5�Zw f���dO��s�I�X�B3�ImK�!�Xլ�̲�p���뒲6�%J�1�:Y�d�9B������µ�AK���E�1=J�"��\J7y��yr�c"�I;��ql�<)�bȴ��n̬�4�,�6m��b,KVh�.�]�Y?�
'�=��:D��Qܡ��%��^���:n��^8��s�UP+�?��+g	�j�|�����ً��g�OB��*�Ґ[>�I?� $AG��%�ooS����� �Ɏ����i��~���L~�,g�}�~]��ʰ��C�ЄM�<(��D�8`��P� ���<~���ۗ��=���|;������߰4��}��F�z��~ΚkYK5�ɕ"U�iM"�\�И��	��xR��u��/r)�)�2���$c�s���΂BLY�/F4)fR��H��5�֣C��=l��j���/R[�x<A�%TI͘��`��B�Q�$�	7���댂J4�kb��K�jx
5�i����,}�~��9�=��6��#ML��Rhç[W���&S���%Jo�8|Q�41D��h
�0*h�X4%b��ʭ�����c_�޿�(a���r�]�"�����␫����=��0�Ѣ@�A�k+�}���Ye���k���#;^�Ο�e� ������FRf���İ"-[[c���^b�Zj��8��w0(z\k����@|���5>��ax�aX0��@9z�U�u�y��\���-�_+�	���b�'?�	�z�)�Q8}�x��֘8��lm�u�5.��i<�ǖ�����,X(5�C�j7��uK��@,�ːeT�m�̉����������k�3y�Ν�ń���R�b�[��`mPB�`�*�|n�Aa��΋��#�vD���|�͸�sXk1�a�CBL�)UU�!��H	��e���#�@$p��߇���ę3��0	���2='4��l��q�~˙�vkqPz��1��j��^�|�e�-�A����ٛ۞C߳7���$��vĘ�Qn�ӧ��V����Сnh�c��!���#��Iy����{zVUӮ�9C�[��_��hJ���Y�4Y4y�
*'�\`]�7��_`��C� ef�z�d�b,�~;d'�̼��F�ޞ���M WU���0�#6�F5q�0}�56�����2���8Gd����gМ;���W_s���a�d�Bj�da��1�G�GBĵ��D�I���u�s�~�8��O��y�+��^p"F��8��ш1�J��Mt�F�R�%h���!0���V9���L��~�oV4j�U#C��RUQ��u�Ua=I��9�� �e�>լ�g��od׼��<�	g��&����HM�Z�C�hH�!�듶���`�`�e��iZ{�b\��0d�:�
�x�V3�:��е�ہs�^!Nj��,�[#M/ e�?8Ti�����(�՘�&�s?�n���}������]�^z���a[�]H1~��r�ubL������MJH-)D�ɥ[��ѭ����29klf�٫{�)�2s���4��{Ϊ�G��ԢZ��4W����!��$�>6H̨tM�+�)��@�`��}�3r�l�b C$5S$Ai=�CE��}�!�D8��x��j8�x��ǆ��ARd����`b"�@%��Ac��j!
�^�f:AC����K��)4Q��I)�è�R�wB�e4��9����;�^~�F����ib��Ν�
~
�i�/b�eJ�M�����8lG#فKV�3]P&֐���`Be�Z������-%e9]R"Ĉ��~Q���Y�6R"���J��J�ZʲG�E�h�SL}�je��{�a���x=����|�W��e���X�,ٚ���lh�=&��n�Pd=j�&���\�����]{vE[q����	$c4��<��#e������v̙WRR��ar���,��	_DrV��1&�w\����̻�����H��:�UOl�ɲ~p�k��a���P�1�P:�)��$��Ḅr���H�27��W���,�e�pi�Q�)�25+���xk)� R�L��\�"����b���D��|���ƈ�@��O2����M�5�� FS��UF�u���R�#H�X�� D�v��p2���6Ё�'ݵ.)Lk倲j�a��-}q��hAC��+���s��\ڙi���oA� FAvs�:5��5�S���oֈ��?$T#F���14�&��ӀOg�0=J_`��0����1�R�w`?�Y��F6Ϝ����c�l&\���X?w�}��,�Ʊ�[?\_��V�(�:�w�[�e͔{Y��]����]Ѭ([��%
�ֶS�ڛ�-�䑪8O�4%��x�g%uk2	��Yi���?;k�{�s�򲱡7�B̓c�����a��U8ek~��{I���`q�P�mf�u�<+.]�U� +e�K��}�+;��������b�¢ڶ�v�;#_Rj����e�G��(,�wH�?��H���F3	���Ā��0mk�$�Q�v(~�{�"��I��y>�6d��v�6{F\(�.[7���:���hj�uM1m��V��A�Ɂ�J�V��ޗ���UH1`�+�ẁ]���w��y���.@
�� �+lv��A��Jh�ʲD�3m 45Q�H�2�� � ji��(�*)��_b_�����Lx��|�C�=����a�k�$�+{lT��Z˅��a�c(?I¤��6D����=���]{����O�Rd[8I�떏�3('���0���K�J�!ߌ�LɎ�Z����TcM�	�,}f��k�g0��|���8����f�����}�Z�Zl���I��%Q�s�C6������]f��f%�e��o�LȎԪϾ�����0d�y�Y�VL�(4���F��"DE��kvX��eq4�J݁ �b����?eF�D&i����2�b���hɍst'�j�F1:��UaN�"F��г�Mb�F[H��������ܻ�%g�]%��`�\��vkʻ��hN@4_��Nj5�C3br�=)���{Y-�@Ԙ�AH�Ċ�����*U�f̉g~��O������t<a�� �Gb�X��0�nc{vx�n>~���J��TT�m`�N>�����_���g�Ѷ����u��ÏbP�c��4��V�?��=+u4��bL�)��N�c="��ڶ�3���0M��%�����y�E�m�)K|P��8���8������Z�^��NH%A)�h ���ER����1���"�y3�@��8��tdge��e��R��{����OU��Z��ٲD�vQ!d�'Kު�h�(	��G�%)�dRޟnG�j#���η�Ϟ���ֻ+!�<�����.(,���X�#�Q�jNWh�D�;k���:�ݮ��ْ�m�S��4�.0�
�)�u�F��*����4���}1���g�瞾�,<c$���#|��<��\�����cN=w�^+��$4u�fo��
{�һb�/��S���8���n��^�}�vlϡ���l͹<��goKI퇶C��>[GuE!	q�9v3ؒy��lQ��d�3Ô�Ѥ+�;�p.�t��o��^/gg�јw�Q���)��&�}�xl�=�\

aZW���q��U|Y@;!u�cI�=�FP�
�v���WvR�K�stڕ�Ӯ׍J���l��{��<��8#;�k��;�YE`��(�y ��9ŷ�A�.B��<��.Y�(B���I����ag����w�T�e�}��b�����/}�t�߲��i�dGa,=�LZCԄh"�����P��(�Sg9�wρ�>��G�[^;��o���W�r���Ȥfay���.�9K��6��w���1��&F�*��,����2ۻ"��{�G`S��t�vh??p����ьڀ�HtB TM3��LQkM�����SB�AR�6�����[7!:G��b�����G������<VLn�jBb�z�z�!�5���˂�5�7�Y*iv�Я3Y�J�aDF����o���;�R3���Ҵt$w�龧�⳾�l�)���c��&d�z�q�h'ʲ+@�{���Z����R&q���۞��QU0�̩J'�#9�6�����0��5�ٚ���j�Jk��wœ�k�.��������e�<M��A���Z�ު���o�?NZY"��f��g^f�����Ø�M��7��}L�78�0'������^���y�U��D������s�{v��zO �#�����1�#���ICIB0��2˥�6�4�-�,)���6J�D$��h�x�xeo�F�$�j�}�l��}wһ�.X\C�D�É�Z�t>����3��3��s��a�����Χ�����5��&
V��u�K+��+)Mtt���v�һO�~�(jR��K���y�S�U����Ŧ;}kɣb��b������s/���VM�9z}�;�����}y�Cs�a�˗�9�]���^�]�cM�	�������!Q�-���}��I�_5���8��D,\w����Yxϵ����7�O0��4�,/2=y������d��7�)��bڭ&P�f/K߳Kl�jس����#���&��I�u�BQ�Y۪�l"h���bQc�d��`3��h�i[����e�1u�ж-*B4B1�h�}�~+f0���_u�k?�1����p�#iv�� :瘧��{�`<���P9�6������?׮�5�F�.yJ�/�a	_�h�(����I�\v"��%�:���i�����Tr�^q�J��
�v�����gc};1�ݕ�fǪ�N��̾@�q�D���BG�v���Q��yRG$��;�K����Yǽ�͐��k|Mw}���G���p9.2���5���#ƒ
�I�4��_xdi�/��ۤXSDe�\�bjYa�o=��;h���<�`k������z��������O�I��ĜR���/�nog��ɶ���ln��S��Z�Z������7'[�U�!t)a�t"&��cS�X��66�����#���Cf��h��\wz�L�����@w%�!H�&=���q��!��v��er2���7��r�_�1v��V[<��?G����^d��1��3 K�ng��`�2�Þ�2w��5����<���2��U���ګ�H
N��	�T39C���9�b2g�I�|�k���e���L�����ສ���0�|�woCv���ڼ��u�f"+�4K�2G�ͷ1����4_Rbם.H~��8hxӱ�	�:���&����1ˋ�d��n9�q��s�9\��ʇ�O��;��>&'�q���-s��腚��qc��p�wlZ}��U�kJҶI(�ȩ����߸���ٻ����p�#ň��	���m��������)�	��g�J-����(�j��x��H3ަ�S��9&1��5��hL���h���;�F�i0.kP�$P0����[>�)���#yK���rmT�7�I1#�mc�M��煿�[�~�qU�eFMC✜�����MJr�]���Wq�m���[�?����
�nG$91i'K�t�-rfmw����Iw��]jjfO�<��GƘg��kf��6�Jx��K��y�9�$H�Vgsު�(�2h/�f3�v�|�tI��bR��z�9����ΘN1OvM	�}���r����O��6��Qr$��O�����V.�LhTM�)˂�/8S�U�����҃��Y=���x����;��'9��������"��E�Z�D'��4�����P^lCb,Y����m��6{��=��g ����!&�Ȱ	տI��g-aW���6�Ǹ|���:*�	&&�(�D�D���-�o�����O(G��'ȁ}`��VL669�,�Yԑ�Q0�O�<g�p��{Y��}H��9 ��L�S�tB�la1B���&������{��ıl��*�w9�]`8�Ӿ�������r��3���̲ڹ��]�<ٟmv��}~g�k�/ݖ��K 3�ň��*��C�܋��E� Y-MS7/�F۝�v$F��R�b?����v��h�f@�7��yݧ/}F�")��a���jL[8k�6MU�/ d ����� �}-`+ �'�$8�162��d\�8u���/F#�J���i[|ȷ�o#���S�u�vπ=��g���}I�i�"�qo���ǖ��p�V\�����Ūt�I ���C���B0�J�@�VH՘-Ə0�!I�bb|q��M���=���8���YP�fxjpj����:��%�~���n�>kM0��DI�|u�"��G�,�i�_��׾̉/�=r�,W�����R�v�i�vi�<�}�n"�73���]a;���<�e��{�2�9���9#�`2�j
�!+��Lu�%�;`�n����1���ݘ&";��3仦Yv.WGv3��
�8����b?��Rʒ���m���y�^I��s`mI��1^��?�{n����ǭ-P�y��/=G�"���0��Ȥe�05��Y���KI����B�f�{^����!��ն���'J�6����m�|�$�i%%ST�nPq#���4�qm��F�i�,Ji��TJ`� -��M���>��M7s����u����x�νz��F=ڪE"X�#&��X��.w�ì���Ƕr�i��c�1�ŋ������W�����&a'l��eV6e�l��{;f�+��ߪS�gۛr�������-F7���gqB��C��8��R�5uSӶmqH���b*��%׻2�H����1�������������o� A�z
)p�X�[
��/K�ͬv��-
��	zX����s����s��z+�lHm������;�=����_�6ޤ쏐�E�',Yo7��n$=�*0mQ��{���ݳw��9�w�]���A#�H1:�{�m�����`<�hCP�&���Y+ݠHF��,4�{V!����$�-���E��n���������D�Ё��~/�|������⌇ �-�l�����ླྀ�k�08����5�m$�sSұ���W8����r�<��[����d8�s��������<��r��%�_a��J ��;w~k���q/���@��K!!Ɩ:4TmE۶�Q�F���o���eug��$R�$�7p�];B;�L7��U`�t-��Z[b o2N�:�5��4Xz�C�m*��1�S�
��F5�l��鹧�+����E��`bJ�(Q��f\���nW&����t��F�Ҥ�
��N>� ����+Ӟ��mϡ���G�����	�x�i��5�߽O��m�uzԈ乥]eJ1�^�ͣb��y� ���
'm��x=7|��z�!�UW�X&MD�ߢ���O<ɹ���D���������u'���
m"B�C
��Sd2�}����/9�O���Ʉ5m)&5Fc�ݢ�1#�:���e�v�ǿ՜�g3q�ݎ=�κ�߷�ܾ{L}V��Έ�4iS"�S�m[���E;�U;c�{�Bg�.��3��@v�򜜇�ʁ�}���\�$Rj�m�0�8�G�9eA�	��l��1hV�KB?��֗�ʓ��>v�B!=���M�3}J������ɋ,���"$��9��sA�M	o,�|������\a���l{�]l�ޓR�kL�
��=ۚ�q$�v�+��Ƭ�Š$�m.Iw�Q�۞u�ȓ�QW�e�3��x�9��C��{���	���a��P��$2t}��G)n����'IbI�����E��^�k AZ!��Ln�0��6�9�~�W���\|�{��7�Eh�n�6#��I$4���%��h'�z�L�X�_�����d˗���"���IS�!G!)U��ĖF#�&�sޱ����R���>g�z�+�Ͽ�ן���Av���Σ��%�Z���E�;�H'��`"���ZB;G�C����Iy~?�-H�Nb��\��E��n)�	�:8�Ҫŭ-150�γ˽��h3����X�ύ�o&�?&h'!�h��Wz�ڞC���@�������/oه1Cc��Y�(�hʴ�IȄ2��͜.��$���KC���p�}�c�C��p)����N ��t�iJ
ia����'~��MFE��F�w����R�=s�NO�L��,���x��+g��m��UMa��Lv0�YC6���n�Z��+$͜����W���?��l\Z�ޕ��.0\�[c�9K1�GY�g{:�mv�f���J�Iq�`�É�W�����ӕ��q4��3���w+��S�x�x7�̮�������c�|4N5�M����D��4���%��5��(�J���h�6)E���ljY�K+L�G�1:t���7��QjKs��/>���&�,sz{�QQ�s��$>f�IE�T�*�_�C�g�����ߥv���@U��p���[����u��t`��jF���.Y7���ώ6Xa��P~���އ���-J#B@�B4�o��Y�Z�л�z���}��ڷ	��w�S��"ͤ����{��"��R�՘ͯ�#ӧ�buc�C�=Mԡ!Hs�t`>f����Y;�K�޹�_�.�|_R��9ٔRfvs���]O�L��<Ș�ږ�s�1F�6���#��~��J��N��L�N�
~Ff��ri�������r�\�הc��a�%�tE��Y�!�fmy�p�a���:��s�?I�A0��x�+ �PR�$
�yB$)�A��r�Mq�M��G���_��=w�W'��8K)�J�p��d\��+���SkؿQ�_W�$e��3�}�[���_ǩ߳� �s��B{����aܶ$�ʁI��E�f)��Й�;gd�n.�W�X�������nn�O=KZX@n6W�ѳ�\&-��v��ڨ�$���>�'�y�3�����G\w-�[�
ޗT㊞/�&�*Ҍ9�����"��,��u��-=�2�M�,�HI�Us�`�Tv	W�D.e$ygدT	���u�ݖR�����F㪢I�$9x����$���d��k���ZK5�RmM ��C��I���3]�7��p��{Ҭ�'"8��7������9��bPRxG�� )m��5��m3w��Xk(�ȁ�&4Yl'w��1���m��p��7��G؜6���}�kVr��n����'�bc�"Ep���L+�����?T��&)	a����ߍ�w�߅�RxBHLCB#�D�������A�d�m���C���9�������^���Eh^}��S�	O����������|��T�Җ>W��n��jkq�3������?�	�܍�F��J�B�J�Np=��L�G^��_�;w��$|[ab���4�Ё�rvi:�S!gx����2�gon"k��5�i&�4I�c�
x�(0��qX��!ޡ
��1�锶��X�tpI�#�Y�`f��.3���!%�*M�ͽ'�&b�v���a�|D.j$ER$H�?�0�e<C  t���g3IRC�������EC_J��O��>N&��:�٨��[Y��~����Wi�W��%��6Ke�1��-k�k���N��˩��з���&�s��2;���c�Iې�V��#�(��w�C�Z�C@� x�ܞ]_9��R�Q|Hبg]�^HA?X.�t��^9��+gX��o��{;��E���5)	b,RWRk�\r���t�m���
�Ct�F�R�(�ح1\�H��'x�/����`�[�/Z7���b̎b�x���E���T������ϲ��}Jw��)El�I��N��n�F՜��|I�o��ٳ�{�)3���0��.'<c�3���h��Q���B�~LYEOl�۞2��hs�[�,����r['��eI��GD��S�&�Ν�&�{G�|��k�T$
�x�e�L��cu�ba������HM���BVV@,Z�������w��6޴���D�3F؈�4D
,���an�����b{�]fkH1c�M�GH�nE���$_�р1~�~	�+Y�ʅ���;A����`���"t}Ud�?�d]�?����]w�8�CԔUќ����ѻ�ZF&k�Ǫ�JV�jԡah��ϟ������y�b�h�xѬ*�Q�*Y�k^I�ӳ�0s��?C�O��n̞�|���m���^���v�69{6��,^2m��<zY��Jq���JoF�!�л��E�[DM;�h���H.�����?����K������_:�8ۛ�:��&��)�9��`0b�Ɏ<�τ�>~�p� N�,�&��(PG�*L�;���d�X>���������<��7���qka�M��4�9E6�������g�<��M_KJ;����x�#ܳw��9�w��~,�ۆ6DcS�n�ԟ����QOl��.;o�:���(ݍ-%�|Q�Qɽgf�`������	Kj�c���S�>�<ͳOp����� �)	`�`0��Z�E&��A�I�\Lѣ0��N���4/�/�/��h�'K>	,h��rf
����,E�9�ԥ�����(�@�4����,x����b/oF~�ڝ#���L����DJ�O���gۙ�ޑ�_��>ˎS'B�+�P�o[l�Ĉ�m�|]D��0*J�a\A.��S���*Q#R8��;IC���"�E�w8$˔�zW�K[���Y�Y��N�~�
뮳�{�^�򫹐��$Mhi�Qe�40�22�=b�����-��*1C4�5e5k8�AcŚ�Ć[�k'i~���,x��y��'x��`{�m| ��d���	��␸�͢I���MѴ_�I�s,��6(�%^��A��������E�ІH#��$�}	�6��)I�ɽs�LAkם[�T'�8���ج�e���� 1@�&�f�d����ᅋ�x�[����i��Kl�G�N<AKIj��Hh�����3<�'����Y�zzI�I����=h��ƈ��U:&����/����I�����{֭ɂ'&�#E*�=���~.e���^M;i����3ʽ���y93w�8�d��q��Zh��4	T(���Οc���]����͔r�$Y�m"������}���$g���c�wZAz٣\�K7a��
3;]�!�2E �|Ik��k��k1���Ʊ~�")&zeI��V�b���S�A�H�w
5��֙��'��ns��g^|�����ǁ?���*'���l�p���ǁ�>�s�7x��@�=���	��D��{��ޙ~��k�}Mʸ�Ѥ���C�m���R�SW�,.dB����vQ�f�l��84�b�ՆV�Om�~������]�o���ݥ\�A�iǑ�+c����P�+�IE��'����j��oN-)մ6W�*����Dk�X���Nw�+��Y�v�����y&>뗗I�13�)�`��ܽ�%(�&
rs�R_>OMg)��c��_�R`�%��)s���L2cL9��)=�W��D?�����^�$���	g,�Y�1���G %�j���������;��ٙ7bf��\�wN,��B�HJ�j:�;GY��<���Q����J��R�g�)��������t{��?}���Go����|��w߃}�Y���΅����9dK�f�i]��7���i��u6��'��)��؇����	���mϡ�K�0B�jSb\	�>U#�]6��F4��A�M�$�l�i����2Ukq"�)�Ք����^���9�'�����~�^d�~(��0j@,q��1��c�������a"Dڶ&�Љ��11d~�[�u�WWM72Ri����=��uf�d~����芪Ep:�Q��٨�1v�yV�� ��d���9�����(2.ߑ�}H!�[�K�Mj 	A�-���[[���kbz���PUĦő�w�(I���db�ԕ�E:H�l<��T�of�eU���]u���Q�8o�{u۠m1����kYZY�����1�a�P�&�	�|   IDAT�����&�@��*�8ܠG_W]s��;p���-��(��g��;)|��������%��.n]���r��ƹ����b^YoR"�D��ǽlϡ���ǲ ˤ�!E+1�y��?�6.������HQ2 N���gы�"�(mκ&	�t`ʹ�����Z2�|���5,=����:,>�ؘ3���~��/}��C7e(�i&��S����2�3����D�G���/�"�5�l�R�]��<0��D�j��{�E4���2米��` �z�~�Yȣ��*v7/�	wL7����g6�)�����#�2iE�gRM1�PxO�"��!�� ��2ٞS�3�)v���&TL��w��ɯW�e�2�̮V��;��H����Q��@]7�R��`��m[��,./1��T�)!4D��J[`��id >=���/�^x����������;9�ɏ0:z5~P��σ���U����]���SK��;�G%MB`�^�e�g�D�s���[�V��4THL#b�dJz�r���9�
�����]��@��]s�=�z'��Z�[�Z
cp�_�8a_a8}�?���ȍ���o�*�0���69;��8���%�3OsC�I��jpi��G+ӡ�Mk��#;�Y�T�#I9�ΩZ�мќ�/��e.)�&;�y}Va���d J��|�>�7�r�t����%9�)~�����C�aq�@���s��i�)1���R8���m�t2f{2����gpF(�Ǚ�����X޺LSd����%N���\b�J�4[��:A�@�|A({��%��V�;<��dBY���*�4-1E�	�pF0�P�ݡ�5�0�����+/1��?g���	�۞�x��ϟdPE��g�W���Ӗ��g/����qz�I铈yV�qn��{�!�}��F{��c{�n�}�1 0M	5N���������&hd��D�]SZ���Bʓ5���ggޕ�ۀ}�l��DE����5�=���?�K��9��o1)�=}I��3��'���W��mI��_Z�����B5ŗ�Z-Kk΀ш�|\��� E@����P�	d��;��B��I��N�_�D��N���	0ٱ�Q�UZ#��&(� 2�t~KU;���%��X:��+_3�6%�x�h��d2�N-�;BX�X�[ˠ�'�@
m�2BR��H1�{}zE��6S�j��et�z�/��kV��K��H�D�PO&��3� )�jJh[b��e��@L��xLY�,-/1O���#!er��,	� T��6@XqF��:�*��4���ֹ���}�&��0*��z�����QLZ֊b�bo���%#�Sb�ȱ?�5��C��Smϡ����O~/0mBJX��F���I7_����s�m��B�1+�� Q�"��d�y��eSƠV��g�����!4�S�e�6EJ����M����g8����ʁ��.-@����9���8�6Y��97m���P8VuB�#��cʒi��@12���hc X�K��N�Q�O���I-�糳1Y_;��:L�� o����Jۻ���L<)s���8��AS�gA�5��<� ���1JBt�mb���$���<1�%%%U5�,/-qak�6�ksY~R�!%�1��� �y�(}��H1�Հ�R����mϯ����o�����NL7{����X;��8r	e��XCU״��t2%i&�q�ዂ~_h�-�&PZOU�xU���Z�q�a]zF(��ԣӆ	r�w<p/eo�+-q|�W~�]z����,0$n]d��ɦu����\R�n�R�a�WzG۞C�JQSK#�:I��cIZ�z[u.'w��
�d�e�iV�)��\�Uc{�,�juȆ�q(|��J�qxW`��9�V&-ה}�g6y�?����}�y�8�����'���P��T����q����f�:$ڢO����������8�&Lő�RB3�W)��e�{%�h��"8g��������b"�X�Т�`��h<�r�$ePdP�JQ�l0�{%��0M�)Ķi�X��|6��Ʀ;AO7oP°�1mj�ؒڐ�eEs���#�����}�I_�J��~%H�?��g��~LG7+������@����k(M������7�䵯�U欷�������6!���o�#�1��ê�$K,��9���S~�P�������2/��_���,�G�d2fuuax����}1�7U��
�NJ/*�?� W�e��H�s��P���>�e���bb<8��u�-(RJf`3j�d2y�$�Q��u�7�<Z��Ն�6�aci��O>��Gooc�>V
�"�?�؞�x�ɳϡc��pP�����o�<�%Q4����;� ��
�����=~���m�����LN��w'!l�Cn���;n!.(Jlh�a��/8��'h��CE��Jj[�E�I�_A���Mh[�,S�����T��4��)�L$�Z���O��D��̎���ywe��WMtH��y�ܗ�U��~5�	TE/#�UhC���$��@��@�rf^���Uf��;���o���X�9��d��V�����ٺt;��Ś<Z��*B۶���Jڪ�"X^Y%����^�oSMk�K�����ɒ��*�%϶���]���0>v�S�c�#����޳�ϾD����P�V�1ݸ �V����bPC��~��x�ڞC��jY�6�H)��`%��K�p�
���QHD�	�,d��ޖ��G�!�a*���n��஻�[B���h�IE�o��.�g�V�C�톋�Np�?����P���ƒ]���ֿ�=�N�ŗ=n��f����>�V=慿�;zKK�����ޛa����]V�^��6t��~�GTM�!��X�r�������Z$y�Y`,�)Z��>�����CW�W1�?nd6ˆ^\���~�k��ʊ(�zJ1�b�/qM�[&h��g%�lWR���?nJ#_P��8KҴˇ*p�����̳������=�JN}�2�(A�6�MuI07�ҽ��Αө�E���*4&�3hRb��5�m���[�[��@L	�kf�$ev����k����0���`<��s,�`�z�F_b����:��t���`8i���I�:�|3a�$¢U�<�0���_e���_��9�w����� ���5111^3��s1���|aʺƚQ1����)I*���.�
��`KH�����!#B�����)'�;ƭ�� �7Q��,����?��4&Z#��,���j����1�E��_$�쐪q�?���j-8t�-.ú/��=�_��2O=�$O|�[�q�Q��6�w�����֋'h^~���ueF�����k@���Ec��8Y�����}wһ��;���?�X��۝���3�3<}��?�	�<�M�?�,+�D�FIp��N��Kb2��
��Kzغ��9[-JK�Q#i6�YV��9�\��%@����N�hd�MiS�N�ih��U'��B�OCa}���;�:��B�YO��^c��L�������jP#41u�p"Inq8�X�ԡƜy����Z���r�u�С�ì_ �B��S��Ge�8s���	���3g[ML�^��N�=�����h;%��� ��'7�}Ⱑ��*j"".g�)f�R7g6�zw��93s�]��D�F��@؈�~�$�}�)z�!��L��m��&r�Λ���� ��z���/q�k_�������)7T~D��n��c\{ۭ�b��=&-�z{�cW�`!y��s�wУ�Z?�Ͽ��|���>ǁiÒ/1���T�L�_�f9����J.	oY����{�檏=�����}����+�y�m6>� �������u׳������s����/���C�8 -��9j���e�o���Ι�v�9��z�5�C�w���gv}��^�|�~5�NU%��2i�T)��;|�3x�m�(^Y�����c���4MCl��'B��TO)�^�Q����jʴm�T��`�`�a�H�`�m�g_�<�?� ���i_xC�·��?�#�f$�tRS�����Ģ[XX�&����o�җ�j;���ڽ,�h{�f?���IU�1Í���^O����fck=����v�8U\L�ݨ�\z�%�9י��{E-��ӬV��C���P�uAQx����{�}���` �4L�
O��Y��6n�������l.����ko:�Շ��mu����0m�k#�~�~�����3��aϒ\���Ɠ?�;~��������o��v�<jy���+��&+E�
uf�����o�2��o�.i6 ��ڵpo���Y��`5�D�u�-zY�ۗ������>�(G?�	��7��F��o=:�=:\���I�aL�CW���_`tõ��7ñ'��H�,i@�R�m|��V�).ſ���ؙ��`.���;���f>��J���.U�]�������I/��ϛ�%���$�:k��il��-I��[,v�;SB�BKT%��ZG
�^���8
�@,U7��e���IM/	֕8���Q#��D�6D�J��(@
�^$�gNs�/�����/�����N��3"����B1*��Sj�>Q������C#O W�&*���B{�����;�VʂUHҡ��o�ꇮ��Lk�/a����T�D��D�ma���&���c�ܼ_*��;��"�qb�:�5=Z����1�z�Vkp-㧏s��ߧ��r�C�b���~����Ͼ�ᛮ����R؇?z#Uy��_��A���EdH�P��[Y���Y.R�=�S��p�p���XZZ�ڏ_���{�y���믜�&I��1�=�9�w�H�Ɩ2U�B9�4�*�Aٵn�.ޥ&ڱ����qy�_"�t�BLɸq�p��Q��������	�ڍڮd�9R#��R���(7�f \��������!?�����+�E�P7&�H2�$��{�v��2��x�5��e6ǎc}t��]p��fX=���Ok�|���z��]G�	�p��IC��('�����X�q!�,S$��BLL�	�����j:E��?`T� ļ��P0�+�*�R]S8���"[�L�	�F�Y�w��QW�0��l=�,[/�&X��$��~){��+�Po������ۛ��8V5�Z��S�*�6	��^���=���W��HR�u ��\�U7��[7�'��S2�+��:�=��{��h$���u��8��m�D��ܚ��	g-g^}�~	��Í���6��=ߧ,@=!μ�*�_>�ha��d�Ho@��c���/Dڍ�����٫�X��}����F�՘�2!w�����W_�O�7X䎇>�{�{�J��~�3O|�����Ba�Gt�:a:ٞ���.ė���yҜmД�0sP��ەf�����K�b+R��IE�4d�(�p��4���gPZ�"����y�<n��W�r���~V���Q���n���/��O�?��*��`���k�|���9Lb����|�q���:�l�.+������{n�YϬ*p�5�6,o*��5iR�z�F��S��p=_��2��S�K&�esk�(�h��S,-rac�`Ѻ9.F1E���"�N��x2�0Rbaa_xD3�t��<����,{`ml��h�E�������3�x��?����+H
�����5ts�"���?������BJ��2����?����c�{'؞CYa��$B��$�yl;�-��RlѪ���s��HN�w��%H���H�찰E�g��zL
$LI�-~��G��y�w?�����G8x�=���'�&�,�bc�,�	k=�C!J��H=ޠX���D�5�5�z��ʂ�G�Q�-&,>�0�~�#���|�{����">���-�!C�hQRWujhb�t2����X��h�7���)��u%�K�I�����sL�!�%E�Xty��Fh��O�⪫���c>��g�ֶ*b2[�L	o�VO!f��I3C�N#B�ʽ�2}�E����S6��"���!f������������p.h��ޅ,�w�o�~�"�8K[��	)ᬣ��w�B=��5����ʞ'�n����0$A��3�����=�����D����
������4�H[�,�9�Q3W@������\ ���J����c�[��|�y����\G�C;��D�{HJ��%�Sg9�[����%����8��U�^�����;����;Ď��o���6�Z����7����A�H�P��-M�7����%�y����׺����I��&N`�<}+�6.���_��b���;0���Z�>x?~�	z�v�?���w;vm��#^<[�8\ZV�ү6	�Xo3��&�moB��˰��:}��v���5ܷ�)�}����ŕE�����p�$k� W���b*�"���R�P�H�n��A�G�\~��yf}ɼ�����٣�2i�&aT0)!)�X��\,���y�C��� �Ec ��+��vɾ�q�0�����/�d�~/X)3�:
1 �K����~�8�?�j)� Mu>�:#��m1�t-e�E1?Fv{G5�������WBǩX�q�!e��2|�p��k}{{̩S�)�%+����ca��
����k�r3�C�1F�)R��*�?�#���E�Ϝe:�PK5��������-�u�3�*L`b���m�&A����z�H����nX�UՔ�)M�6,������L��im���2B�b���&!�d�S<̡���o��9�w����Ɗж�6L��4�ϥ��+�1�).	eQ"1�RBB �g��=u���Un�Щq���	�Z|3F��B��r�&ַ�8�w_�����]�ٜr�{��k_}�Ϳ�*��1���Ρ�[���"����?rx���ѓ��U�P�oR7/��Я7���5�79Z'��!�Z8��'�K�82X W3��^�����t��m�8�f2!��8�tT��9�Y�]c�m�L�j5���E����7���J��A�]�8�P���n� Up����w����<��F`���fh�"�5���LF�@�ٻ�	�8W��=�����e�c��cl�?A��20�K��=�<97]c{׻.�л?�,�|۵f���#���*�:B7O!��ټpF,I`#LEa_�ib 45EQ�I���b��ŉ!��F�\X�W����:ަP�W�U�q�6tD>@�+�EA�Y���{K�=��0Z�e���Y����o��G��{�®�Ro������w����9X%F���Ȱ,���y_��zXo�Ҵ�����Wv��%lϡ�l�(P�)@
^b���6~l��#.e�u���6Xg��p�Sg���ewC����$ؤ���:�k���_��z�7*��g�������Z�,l+﫠�O?d�?�Y(Е�����.V\w���y��βu��h�Gz�y����\8�
'��OвO��q�o���������ӯ��~z�`�0o���7α�b��&��$�8J��!�s�*���S�J�uv�e�w5&��uNk6����tI29o�&j�&L�٤X1�+ز��b��?Dq�uhѣj�Y���&�DgL��Qu6oMk���fV�ɂ6�:l�ud���2~�ǜ��k\_�H��[>u޻�E%�h�[�4G��|d�z��E4(eW)�F:\���}��^���qP7�P ���"X�+|n)t��8B�`���fc�2�%A��u����}pz�,�V��Y__��*����g-�HR�� ���DL���ӆ�b6Οz��ʈ����?�<��5�e�Y��v������������9Ķ�,mV�O,��T�wA�$�,g|�����\�=��d{�7�~��OcE����	")���>"7.��Wc�X��U'I�M^Q�;*V3ёn�j7"��JSj�t`&lG�L�~�3"B�� %�5�o?�)SR�>�p��\K�+��0�H�"K�a�)IQ�Nn�/D�U�-��O�e��y�1hY3�U�fk��ON�B[����&�����O�Qj����ň�pB
��6M�Q|��R�(����;��,K���!��uk�]0%�b�2�5��zZѳ}�u�����O|��{!���"b�!䊀Es��:�؝���[<j'�麖�5ؾ�Q�ϒD�������?c��q�x�X ����Hg�4�!�w��JWb���͉Z�u�]�3�Ν�\"uW	?���k��.�^�K.�ˮ��p�6D
�IQѐdڦ!�@�
ڶA�������64gIuMմ�����:ɗ��5d��\��B�[C�W�b�5c�Ĭ�/F��K�r��	
Cj���˚����\��㧎�q���p#�y�|��l��iʶ�ޞ������:�X{&�;ۦz̻�bݹ6F�6P������ٿz�s��Z������1��XٴTVL���p�Z�1�4�$���)v�P'�;�z�Li�NA�� ���M7�]�H/F\�|��Z��gb}I��"�"���%�Qz���&bS�����ore g�bbE3�NS�Lc�h�R#�E	�Ä��ť�ilKh����RG�,Y\XĈ�yO�ִҲ�[&��d{���h���n��:O�톏�c�����Xux㨵E[�\�-�M���[��]s��+i�d� !ktw\��cJ)��������Ir���ۿRv����#0��z=� ����R�D�-�$��w}q�9�3�6ف��:�\A2��w�
+�JH1c���}ʏ�� 
��`�|���9�_f�� U��Ƕ�F�ŠL&c\�<��<�VWIF����4&B]Q@2NktR�bB�f��<q��ec��9@�,#L�S�&Z���E��bg�7�0�V��R�iʂ.��^����O?�~��o����￙b��a�Lq�45��}Z�Esa���������9��&�j�BK�<g|��{Y�o��9��`��oAi�B��MU�ak�G���f��@>�Dh5�RDcĤ|�eK3���6<cǚeIo&��c�.S�,zi�I�BB¦���)��CFY��K.;3��"*à\���2q:���L�b�H/	���`��#�-n"��D �0(A�T\�a훂�ވ�ﱾ����wXg��7�s�Ϝ"4-�=FM�;4��q�:��l"�b�"ML����̸����Cq��h�#	x���^tu?�
�"�Y��{R��w>gs��̡Ana���|��?x��/<͚x$��Xb��l_l��K�E:'{�����	!Zhb��@[U󂐈��uŪ�t�~&��ߗv���j$(L��Y\\b{�ͤ�R�J�IE���Xz�g0������	���ڻ&���	X�I	3���i�!�9ۍLQ`��z�x2%6M���f��[��R#��$�P*W3n���/�Z����	������>K�us�fͮ Z�\��b�L��+�y���>WX}REN5	&mdX����{�����q�m��$M�!a��lL��j�FM3X0kZT[4E"�ZS�c�$�LCMZ�����Lla�X�i+;Y�_���R��'Y$�*�
8���/dmMP5���&Q���؄M�2(��K�6��t�FI�K�>m���i�Ր��11�b���VSx,�6�i"[^�����<�T5�8v�jZQ�}�7�h��^�O����*Y
$�J\ڕ�S��Q��.�ܼ
���`r�k0`SWra�{�鳟��?@J���_z3c��Y�{)�0":�����	���B&R���^��M�X��k�������ZA˂�(U
�z��̏'O���,������5�V5��d��j�v[�]WlUS��)�mŤ��چISq��4�G�޶����1(�MUc1�6��жy�����kb���U��5����?�x�M�]ORR8�XX^%^�b��b�F��HS�LmE!-�?~���g-y>t��?�s��O��O~�$UQp��؜���0Z�US�G�SQ?��|@E�"LBB4#���7��2��P��ogd�ƴ�6���6�o/�?tP�Pm�j���1�	j�$�$�$�$�JJ�<�%j<N�� �3
�7��0��K�v~3�������MΎTD�j�
���#�F0U��� T�4��4t��Y�ӯ�Hr��,`c���ek�۞t�6�='��8�U�SO�˞b9q��{F�+�i�#��KW�E�H�	g�`i����2�y�:s~ݲ%�ح�U!�,�9���ӟf��ۃ N��m
��� ]�j2�a�Ǫ�$�lm��SO3-p��[�a�� c^�A�@���ezY��C��}�O���YB����ES��W���	n������j"�$�زYO����Y��zY�,�L�bb��5x���S72geW��m��4�[,�8�8y����y�дe�����PɎYl����hb19���@�U����Ũ8����r[�+�䊻�c��`�VQ��$��}���'��/�\s���[�J�]��C������_�G�W�q(
e��P�;E�p"�<:�~��s*��U�,����o�흹�P[)T#����p�{�{|a�-�XMD|��@�%$��P�K�)&4(��8�DEb��1fW�u���vw�Ze2j[f���=��AD,bJD
�m\�l;�^5�p����\G	���J4�E[L|gfCx)�p�S�{��Z����*.�11�Z�O�J[ς:�l��%Lk��-$%�i	��Q�F�:<IɌl��]Yy�Hj�N�{���Pԉ�?`�?�������Bo@U'��M�Z�m/h�R�s+9K6�S��/���/���F������Uw���*Ƃ��� �c��A�x��s���q���3�ؠ7�B��. t���:Ooh���'M�V;e��c��q�hF�[#�l��bdZ7�
��A��<r�v�Ä,چ�j�,..r��鮅`I1�b��-
���X���`�Š֐B�tm�����w����c��Z���f׬!�P��aLVIeB��� �c�R`N��ݪ��	��[�8����w\s�N���8��P�-��!fyD����aqv���Յ} տ�c�h4��Q־�OosE��_���o�=�{�EP�u�I*N���M�;���i�4�.$=G[BߢOQx#���)�ք��ҶI-�60
o�Z��(��9h��ݤrJ��"s�WL���K��Z�7h����a{�����=fT��߬:St���2b���J�¬9�ZEm�����j�Ǚ{�>�ǈ�L�a0�����h˵����mJ�1Ơc�q�!�S���t\�v��.)���|vR�`m�I`h<�*�(VV���C,�p=��2���إ�՜�FQ	͕��0ΡM��O=ŋ�?���?u�k1�Շ���Fm��o����G�}�)�}�;,�2����{�s�5��D3fa~��ͧ�\V'���L��d;�;�^YR��D��5�R�ԍ���"e�A�C"yZC�◪�)��FQ�^ISWH���G����7�XT�6FB���e`��y7g\�|V8��fww>��Y�y*$Į=�3~ٽs�Ǎ*� ����"���6H�g�i=��o��u���xa�ko���I���9��Ә��X�66Eh�#��?Z����X��� ����s���o��9��@�YK��:F���O��<�Zoۆd�6����>�������w��	�j�	�4���S��7,mְ(Dq1bR��+��U��$�s����f%�:���v>>����{�H�"�m8"�����ZS�^{�c ��Ɯ�͵�g=y�z�̨�!"��v��e�;ٻ�Q�,=6�SZ�l�\^.z8�8��9��4�!�Ė���7���4�r�8�,�M��E�+�v��X�I��J QR��형>���<JZ]�uy]��q1C�6bD2��Z����/!"mD�[o��7�|3�9�pӮ�n\���[ ��-���~��9L|�N��*ó�\m���B�:Ck3�˩"����m.�7�͕�45�)BYf�����Zl�ђ5�]Yp�� χ�n�͊%�܏N�C�;N��	�y��G�ZQgm�tZQ��r��X�Pxb�IΡ���E��{Fe�Q���$��:�@+tYr��`�$A3�"._��J��h�%I�2�Ia0\�xc�`0I�u@�E/,�r�������?�3������X��>��u^=����~�p�c�>eMLq!��� ��tҤH�,�=���8�s�a���&mKHj����������T�L��am�u�z8`���9r��	T&��N�X?�����Au�������.�.n�܄Ę~zZ5��1_P�ʊ]����&sZ�y{wi�ɻ\�^��^Y!�-e�4g��,��.C�����K������<X��������`�G��(��Ʃ"mW�m��8�۶%�-M�R�&W�ͬrƐH`b^���e���d��q��S?������-g9���"w~�#�C�������O@� �;~K֣7�
E�[8��c:r���}9z1��+���.- v��<�֕�E����}d����7_a-��܌W6�6g�����iv�w���u�ϥ���U(�*x��	��$�5j�t�cb�g�n�~o:b�b/vcwbbc���Dk�G�)i(Q�A�"Hxo��J��s����=_fI����U"3?{���y����ԅޘ���"@�c$��5hM9�c]�0d��[�ɔAG�ԆAȲ�e��ϳ���PI_}4�-ژ<'ؚ���䲘��4�g���7�T�>zlm��&�����;FKCʪZ�L�)o���_z���|��_���J�]��@L&̋U/�;Ȇ���1z�ʒ��xmصs7^L��f�����8�udXU�除ao�_X��ZO�D�B�9������
��W&�$�_�0JPyG�<*����ɑַm��qeI��rܕT����g���֖.⣢V��ʺD�N�i���m��xa��g(��VG�*�L��Y�KT���AhQ���c=.��M��4��0��Z��,� ˈ1�C�O����2�̈!�D�҉^�}�(Ce�:D�8�!L��m��Zh�]'	$4��!�O�.�>��!D�"dI�-�X֊7C�����ۮ�v��U��R����y����M�'�*Ǘ%��[���R% ���2र�tΡi��� ��Ls���x���8�cd�"BD��L]9q�c\L��ȚnG]שʖ�"�h��(��DX��R05?�����Y�ј� �H�>13��J��ׇؔX'�rT�P3Ә�Z���|�i@lF�gF)�e���*>8d�HD��H��!xߋ&�	������,��+�6�Q��~pY��3�p�����:�ԧ	
2���M}�S�)�-i���`H̔9���32r"ƸT����J��+Whk�Bq�>!з5�{%��,���0[�>bc䢊�l��K����]�][�b5Do�� �9�rn8�Vq����bU+��S����G�zÝ3�v3V�`-X��+���l�R�H	j�@A(�~�J$��HHI�Ʉ$4\��9�kf�͢���!Q�?Oh��.��u:�1غ�ǀ�� ����L'DzH����L��	�)6��I��e$����	A��*Ft -Q��`#���\��/��{	��A�@M2Ui�^B�$�R��L>���	�
!H�����Q��Q��vr�Ϟ���LSR7�'n�� {��S�d���S���`Q�A��	x��L��&.͐ez�(_B��"�Z$F����K������[�Кn�Cp�#R��ێa=����6].i�Q�t�I��:�ꚪ�q�'���͆US-2c�ʊ�hD�������e��u�w_����c����Ӵ&���4&�61�0:���(�ex�(��M�^�ԴMΜg���/��˚��U�e��T��"��m:c.kmY�����"F�ނ�������֕��Ǖ
�W(��՞X�+g?SFn;$��HX�,�e��{��ħy��7��8y��Y��٭33��Ucƾbe�GVC:�Ző}(��ΙEęE�o�be�4ZӔ����zbLI�)P�7Z◿�ԂiV.eC��i��w�d���>U�.�/*��[�P���9İ���E�s���������֦�n�ԉ��!U�����XM��\7�д�u��κ�}�X+���/ӽ� ���ID푮�QS��x�Z�E�J��K�PO-ަ���D�B �^m���F�87 |����oD��y�/��c��̾Bӱ�lT� ����wO��d�����l:3Z'dwHԳ��t�22��d&CI�Đ �d�ȳ�a�)�:�r�u���J�����������>��I{]J�֚,3x��X�PRB�i�|]*5��l���B�d����'u�1$?�@��дU�M�>B���5��}�����[�#g��x����0�iS�-����2�V�-St���+k�(2}n
��U���b���J��+W��H���DƵE����w\
33�Z.�y`/>�I늣/�k�p8f�s���^����9Jk���p�8'��J��)l�gO��Σ��n3ߛa9˹tv��S�m������U��Љ�d��nJ!dӢ͌V6���e@�Z��"�-oB+SR��.��j�(L�{2��� �"�s�,C4R���A
"ߠ��!��\��M�`@Tj�,\�av�u?�%&
p!U�|6�*N@��*�Cb%���dni�h@X$-s�u6��F50JB�Qbv���g�S��_��Ș��`ҒI��!4F@R6Jk%���ɲ,�������s�U�R�5�;\��yV�WRG%F|HH�SŌ��b`�8���ʤ�qUSU6D�JI1"@I�Vcu]3�p�!b����N��.
��I�=L�M�絁���D�犘:,_h>kR��0	�c%ֆC���ڈwܫ��.;n��k{���,��?���%�'3P�tQ�>ݺb{�u�b��s�~ã�����)B��{���<���+�K�+	�W ^��dRPV�y�s�e���x�A�����Yi�����>x�c�����jW��e����΃��G����cߡ{��a��qN��
'���pm�(h�F���{�1�㥯~�9�,>�BY��HՂx�S!��!h������N�*�I�.-����G1C���!��q���d<Йo�}�N\U���>}�V�E���I� $%�дye�O��R@�H����Ut(�a(r��N�~�1Z��̉UL�+�lI���J��}��1N���+RJB3��tn�G*��neI��K�B2&��=J�TS6na8��=��d�637�ʶ[og�{?`K&�����l�1�������<�_!Ҵ�����f��1ENf�4��-ոL�vB�I v'6�sb36h��E�zGYU�mM�-Ze�
Z�!��yϸ��$y���բ��R X�	��C_�����X�ƘX!4򸤤��H:2�H W��3�((�@�p���8��Oһ���@���na��;��m+��@wn����N\�v���*�gCTK6D���W$a�JB���<#GU�(�
���=�Gf�TiQ�1ւQ����U;,�A2�u'{bfn;Re���Q�&3T"&�u�^��,.-2^Y�����/�s͑�̟;¹���[�T<m�'�T�_�2��h�<���/���W$��GR�~U�����'6�P6̸�wZk�S�cJ�333y��-1�� S�u]������b@4�#AH�Lv�"F���z<$o���BwsV]����ӹ�F�L-�J��%��utı�-rX�tF4y�a@E���*�"QMh�|�f@}��`mRgk���(���4&��<a ��|�.�|�Q�=��;��d9�"���q>u-�&
�w�c�CX����n�!�6u!����� �,eUQ�5���D!hEcO
�&'�	r}2F����9�uM�j<G�y�2�v��V�j<f<|2|�M����i�����Km�8~��r}��`���>4:16� �D�D)�To
��dQa*����z�1�z/�.���Kg�l����nb���&������;T��N;#�92����3�B�� ��B$��5�Br���X�"6�+	�c/|�sH�Dx/���cks:��UE��
-:|��<��J��ڳ����!DF��$ޥ��҆�k3[v�o�aN�����h�����`�n���5�y����kK��v;��F3A|'j��W��M��>-�1�c�lwZ����r"�)�s��O��*`^��K�,�]�����-�SL�edZ�[-��*���Gd#��d2��2-�>z��1Z�XP�*k9_G.m��5�܃ػ2I=1$QP��2�l��K����~��ݻ���O�۱�,>�W�(�Q$޴�Q�Ԇ�t� �,`if�J"\�(���!�n���o�%i۠Z��Һ���~/���e&WΒ�Ɉ �Bh*f����mpҦ�(
�<'�,�ֿ#`���h��ɔ�(�V:��5c��|mNꆫ��8�(�����ή�����5�� ��HE++(��s'�0�k����Rv������I/�2(��s���KG�����x��������P�)̞�,=ʜK�1J0-K.�v"����9"�:FF��Q�J��cW��<�2C5u]�\Ȥ����b7*�U^h����U{�袭e���2-:��n�@��ѪO���u�#R�fh�1(��e������Vl;��]�@~n����6�-1���r��M��������r���!�"�Lj[6-�	0:
�}��K��:U	ιD)�)%�V��v���h�i��6maE����#��H�$h���&�4���d}�@H��K>P+�RKq�s���w;B�Q��"!zB��<���߯x����o}�+(�-���'Q�"Ā
`���Ј�D��i��&ſ���$)W"Z(|m	>���S��"I˂@zM���=��� �^x�㯼��VY��P
a�w����5.$J���5P�۴�<U�eɨ�oL���x�1Ք"zOf2ZYN�4��.���O�u\��������z�D�Xk�T��%%�Yƣq��7��s��rrm�n}��;2����)�E�����F��A�Id�!��8�p�K�}��ڒ�;o��<ƎoC�S�Y��M���ګ���Vi�v�DZ�\^��'v���^�-n�=��]i���
m�co}��"uY!\�۫Fu���*۵�{�����3v����������eñ��P�T@�'~tH��%�%���Z�ՕU��*��v��օ��;-F��-����K<`%J�u�p�et�mz�.�V K@���uj뺄/�T &��L�d��"ݛ٥H��	�I/� �{v]��=�����s�<�wC� �Mm���U�/-��	�E8��#^d�*��`��{���/~�)c��M;�GO-��1��K���<p��Vז��D�H�D�*԰�e#����>n�O���V�@�P.�y������3'_�4Fd%$RFlm�RA�������}��E�Z�`(^%J�U����V�1����/��$o�(:m���hD8�z��ۏV�L#�j�����ȍI�I��vR��iQ�_}\��U��Ƃ�����z����񘲮�$�q,�V^��l�{���~�����F7�2繟��ҍ/�,N��X�nA$�0��,�r�-�q��~�k��Z�}�.�0}�����#j�3=��Y��BG��a'1
c[#��y�����+��Ǖ
�c�RDg	�Ey߉�>8��;v�ܘ�&zK(2*Y�G����	E$�d,�}F��[h"�=D�T��'�/ۻ�D�bee��`H[Ȅ���ז��(T͋�=�v+i	���"��RV�p)6�O"B�Aw;�TTe���@Y��v�Bo �ӿ4U�/�K�N7�|�qX�ku�CFUMa��R�hmj�J��S@ar�<!܃T��\*l�Y��|���G~�m;���*GT5�,���@jAYWd���s:���ӟ�\�go;��oAt;0J~��h�Kˌ��=3MV� 'Q����@gX����S��._��f��e�����r���ڧ��Z)|��.�w�ɖgne���3CK*j暑c\Y*g��XH2m�L��u�p<Jsp��ٽ�t�H�>�9:y�t�hD�[�Q�F�=��}�X��S�	� )�v@�y��*��Tu�F>*%m�$��ȵA��KR��<�{@�R���/2y���K� ؔǓ+[�ڕ��Ji�Sg�?�ڹ�z���]E�@����zs�YT�1�)ff�Hy̎�Tq�<�%�'��$�U1m0�̕��q�+g�c/~�s�����e��l���.k!1ڴ0B`�c�c'��r����x�<'O��#S)q�&3:�u�:�}�?-`ee�3gO�EH �*�)�Nwٲ�ś�Kd��T5�Q1�!���Рn'��N�C�h#[�#6\L�n��#dJ'T�l4��IA4i���4�'X��I�:)�=�c�R�K����U������]��[��zD)E�ݦ�gLj�#QQ |���Ӧ���Vέ7���U��K�!������DL�hY!D����f~��=����&�%R	��2o��Y^���!bd߁l���)Z��-[�t��T�EOg�ǎ�;8���s[����BS���(�L�*J*�'m�D�o��#���/3����>�w�G�d^cLj��󜢩z뺦��ȌJ�6�4���R��hTsJ�'�<$�h�׺��H��y*['�Y�%i��(ZE�Ҋ�x�p8��k����W�٤ J6#*�f�;V&'�/����D)�=U�_���~�	�M��QQ�}�L���<��?�V[s�ڶ�7��������ϳ[w�T�_�!#��꘢���zװ|j&��'���X�ȼ2K�xƕ��1����mEYV�[¹���YINcN!�A�H[bY2�*.��"���K�3�:-N��;�L�Ou��u�"]2��5���%���2���Z��D�*�E�v�;TE�E�Xiu�k�P��k�n�S��d>�}�*dJ.���v1��1#k�gsF�5��/�M�V�h�$0�RA��m�&J��ϸt'��z��5zPS�x�2"������g��P����P�ٹi<��@��Ǖb	��kr
�BGݬ�p$�8'k�
�u�֎]��s�]�-�Bpd*�� "ҋ������Iq.��ٙ�"��va`4�{��x�+N��3%o���]�iT���C����V�Ç ��\R��x�1n��.��!j�
*�LB������ՅB�z�܆��z�{�8*�bi	"����I$&˘jwPQP���$�U��3)I���`��#u����t�ܜ�F�����YJ_QGJ$�z���:�tF�W��	�gTr?��RdJ%W����z6U�^�My|�P��~���d�(&���}1ͨI����2q���()����\���@@��D��97!�j�`�c.,]`�gnd�c���{�|���~��GO3]�	��j�Q���-�a��bG�����^��� O"E9v�Bz�̕Y��1�$�a���'D�������u�8/�mEm�2�;i!0�A�Ό�S�������3��gue	����W�,lAu�L�ne��݈�3�p���Q��Ο"�u`��("J�P#�8}�6��O��������8v���UKfggWk�jH/��Q"�$(�:-dݜ�Ӣ庨����;Ui	�O��"�MZ䁉�%""T��=���fòt���s��� |� ޑeS��yTP��Ha�J�����P;4��tLN�Az�����'atR��9m��u�dg)^8B�p"����%]��
��w��[��B��*?�������r8�l��N]2%kf.]��_bul��&�_A]w���|s�jd0�� ��Jbg�
/#Y�aDH��Q m�Ib�B�G�f���_���f��Ev�hK��f1$�8m��Rh|UQ�J����J؋̤�Qm$�[sV�1���f�.erb���tuh�V�@I��dFAت���u@��"W*��B#��!yS����6S,?`>�;�\v�ϲnD�^�O�#Q����9x���4�4�J4D�砪�2_dl�f���w8���Q>�<[c�S��C�s9�5-����"|U��3V�Z��c��c�9f����c\I�Ø�2��	I���쥪�{!k+�X'{�Hڧ{��t3���8��oq���+�Ob�d��K���B�T�Lޡ@��@�K���h�Z���Mٳ\��X!ѕg����-v����ï���%�~�?�O���)FZ2�6�e�XU��d>
"QZڡf���vg�3f8�EMI���z02J�H3hѨ�� ����h�O�m�&0�6���}�����3dHI�����J�N	=yt'J�Rj��n��S�q2I�Dz�ARzϨ�S���և�Cm��Pә��z�l��4̤uA;c��+�}㻼��_ㆼ��`��ZR8�L[��C���P�\|�%��g�O�fǽ�ӽ�>Ԗ-`��I*����A$��j�r!6nR����cǵ7p��YFFb| �C�H԰���D�U��X;T�\7J�*&�b�k]v����$� ".�d\dmR��ILGHI�h��s��Vשͮ2d��0F�g9F���� & �w�����/L>�{��O���Z���zE~r���:g��i�菙q E���P ��e��z�t+g��㷎3]��7m��	1�P�|�K����{���͕�q%���ؗ?����x��^��_��/�f��̇F^39-y�l���K�̰��������d���d��ĻB S���>���6Sy�kL&��5Up�Zc����������%f��Β���+�Μb��������6.��<G���x�����c��>u��F��{T=�3�v�"/Սԧ�d:��7�kuPJ#CHt!H<[��g�fKW�>��d&�P�	I��A������$5��}IHw�5!Dr�i�ZIs�%jV��"R(�WegE���{�a,M.n؎��L�j"���6��8��Ƽ��o����:��2���鶀��W3r-�hC+
������s'ϳ��J���W�����ǝ2w��榊x� ����d�G}��W^��˯�?3����ڝ6R)ƣ��UlYSh�~3cPZ��F5���FVL��4+�H�<C[���D�SB���(C�(J������щ�wo2CaZ7b>�u�� ��O�I�N��� �����]��m8B��F#��D��p��5��ݷ1u�U�Nb-M_F���g��Ǐ��+��12�-���֬OF����G�d�2K��ŕ��1�L
lU�E�������Z���1!�]"{	䭜 ��l�K�+��ߢ��ﾞ��[9��VX��[�6q�q����HE�*�JM. xʳ���8�Li�ޙ���*���_�p�47<�đ��aǧ�{�KO~���?��>���.�?��2��(��5C;"�2�2==MЧ?6��- ��ݤ���ȇ�������"%��&�	���F�ϒӚ��?:�\�iR�32m�̰^bG!�B��ɌUc���fn�Wl�('PFCh�ٚ����u~��� ��W�+���o��h��6�m��-���6P�j��4�L�a���~�+��1[��9��V|5&�!��S!#뻩��aPY�ܿ�v������~x����p�G[&�r8`<"b �R2�J���(�(a!q�/�M�-ن����D𑑫X�FI?@HT�[7�1w���JU�mx�Rjd�YA��5�y	�9a9��>�=�d��7U�1M�EMZ�L�"��\�lE�=R$�ng��;oF�p�4!�� �D�������*nUPooS�,3ݚ�����Y-UQ��j�Вy}���q�+	�c���y�������]�\�O���^g\�}S��$6b���� �9�r�<giu̹��6+����C�2�i3����qrD�7�c
�sT՘AY"�G�@�B�;�3X��?vyq�V���p�ԁ|���:�W���^s�K�3u�zz;Y;x�����<������
��X1p��,���dR�GH!1RRٚ�Θ�v�:���㨯�T���wO��e���]Jc$��iC�! e��R�� S�L�f� <��j�"*����f�������l�F�M:�K�&(�I�]I�M�L�m��t2�薤���c����LA�^8���ŕ���T��%��}���9��oPu%���,�;�އ�X�F�8٬�4�5��ב��7��O=�����{�;��"V#F�1�� gk�̠���V
�LF�NE�M`n6��!���hP�������& �"Fir��2R�qɨ*�ޭ��()i����͇K�H���������ukU1�Q���.�Qt	��R�"Y�����_�|f
����sF5�vd��"��!9�y"SS]�׌Ugf���3>~;
�jDƑ�dBr�����w?�#t%~����?&��G��V�yT�s��%�_JW6�P�A��$�!:3�QI��A�Ǩ�$S0:.�q�o���q�j��z[w�6�K�!Ke��8�G""�C��A�F@�ĕ5��g��-3�$��,V#�>x#W�l=��7���'�
�Gnd�������ԯ�ű��k/�IXKb(R�h�x�֒��v�C����������b��9���hr��Q�?#&���M��	�V���c�C�$]'~�y1b�FK�Lf�� K�x *�Tt�R�C���\{-޴�B]�i�Ě�S�3�o|��ؐ�M����O�1/Ԑ�q�-�Yz"`�($F��J��I��R��LE�x�����?�raΕr��D���I�M
f��g�i���(��vs��GX:v���9��i�S\L��S�>;VQ663�{lb=����+�mj򫯽K�;����$3�<ϩ���pLY��L���%�kw��O�0RҾ9 �����b��|����s=��?���4��I���Dh�t�+/���G��Bhb9F(��,�!��������8��m���ڭ=-?�c<b�;"��J��q�+	�c�YF��,��<z{�>;����*���\#%�+��hT�QZ���EH/��W�9�'x��2�n����ck��q�J	�щ#�#^WTq�x�g����[GQ��8 zt�H���17���Ň@gj���)V/-�U̇���Y��*��to��k���o}��Ͽě/>O��l�:R0��n�%)�Nw�bT�X��%�*!�e�v�_�M
s�5�'������5��?�T�W8)4Y�ܵ�0��J�a����O�'����j��)�];8�[_��yT0��!
��@�d�ѐ+�'��w��\C�e�i2�<��w�O��^\���;�xQBJ��
�7P��-�r�>�vL��E��o�m��~9=K�UtrE'�d"(Q	�u��8�`[n��������oX�_�,m�Z�-��Nr�D4��L�t��d5���"��n!)���2�B��Y)$Y���Zh���c���{�,K*uZEN��I�<6R�1"Br~���m\L���M،���@�Ϳ��D�1$�^'��lH;�@��fC����!��������Ӵ*	2u�r8�	B���U�i $��!�0�E�#�1��ڥU�3D]b��l�������y�}:J��cƅb�
@�W�� ^��g�1`]��VH�w����ó&�a< j�ER9KT�8�cj\�d�m���5:*�(Ʉ$��Jbj��`G#�V^`�d��������!S,��%G��P_8G�|���eĥU�Q�*��3�=����ͷ���;5��w���{��9���<����={�s�w3uh������wx�k�ʳ�r��)VW�X���S3X2�k(IY�n�o��t���HcN���C[b�z2ż|����סL�� c4�o�YJk��-wގٹZS�A��RwB!� ��D�\4e��-����(77s��q���3p�<3J!��6�Q�h|e`�М�2����YdU�-���st�Ǿ�M��g�;Q��*F���������HU���"��5�n����x�o��sG��1��~�l�ǴVD�P��0�/?��5�F H^�A$�w�gn�o~�*Z#�?};o!��V�zT�c���ht��t2v�q2��{^'���Yd�M�t���c��L���~���{g߃Q ���@�$�L$�d£�M,!�Z�$*.R�wlg�Mw0w���'x��ߦ']�5;E���R�rn�l��A���hE��0d�ȣv%> �$�A̚�x6�J�.��޽:�Yh�������2�[&��b&�Y���Q��<U�e�񠂢���L��������*��NA� ���D ȵ�Wж�#�Ev_{#��w�w�~�����}'um���;���:����!�1Ey�<�o���JI�v��O^�w��z�A�9��G���s<�G�>��<�t�Y&��P�FD�F!eC�1��cDx����Vn�E�i�O~�L�6f�tbqY"�<G�HNv�ք&߿����D�̂Γ^�O�B��<��Kɺ�� �jJ�D�%�d��$��#^X��	5kB�Uc�-:⃧�jщ�K�����e�����D��T�J���+/�˒W���ܴ�*���1`Z
�6��P�tL�صL�;�NJ,�ڿ���?�\�M�E
%�u��Ϧ"���xu��<�y�@��5������� �2�,��F�媭RE&�LZ&G*Ep>���!AoO�\��o�N�퓄��.%xI�b�Z���ccο�	�8/$as���x�F�1zO�9�X&0��f������A:�܌��C���^y������2=Ũ�H�۞.c�p����S���u��}���Wf�̸��?!�mE���m�}��vo/�Bf�ќ,c��0�c�k�L�����Į-p�}�H��b1�u��nTTcO�gti�gtHF��誈�+%�<� ~󷑋c�Ϝ����=v�w�+�?�H��/s���e���79{��y���+�N�g_��gx��������9v>p���?慵۵f���)� ?�t��_�$���ç���\ޜ���GL���96�����=��"�R`�����̰��;0���?z�u�%�y���l"\RH#Blڰ*Wxg��c�������`JK���s�	u���3���[?w�0����c��]��Fn8��EFo��+�W�u�,�U��i�Ui�~���~���tɷ-4IHl>,)QR��,�*�Ρ�f�'�ŧ����U�3�Q��J�� �/�D�m� �Ti��J;����5e]RZK�ƸEb��������i� E��IE��;���{���}:�`!�/��H�z/�	E�AއF
��P;�w2Ħgk$�U���R4�O"c@FA%$KHF�3�f��7ӻ�6Ԟ��2��"��㚛�a����G5QL;����\��.��I�y1F���A+���6���ĕ��K�����UY�������>�����xL@pf4D]����fz���p	�i1�j!ʚ�eg��?s��:���	�ТƖ�H�P6�5�L�c+�*��2�4�c�\s+Yg1��_���fwm��`�y���%G��ʳ��k{�{�A2���Z����^~�-m�����?̑�W���9��o�r�('�����'s����@�Ϙd�� �����F����J6���F3͏6�|�>���29�.��-�o���;o�v�*�Ա�"��@�V����Fp�PV�?y
!���K2��
Y�P����OmAD�f�+�P��ш�W������&��bv�b��P�E�m�a���N�h;��������+�^s��i�[�Dn`	1��EApu�9�(���亇浿��!��h#k�!	��"!ٛ�R Y�Z�����1�ht�ϔ&�����uIݘ�H�*Q[&� Q!Ѹ��?5Wǫ�5�� E����C��w����u�^&_�����u)�AD�8$N�Nq�Zo�Aj �BD:I��Ri��l�ԃ��ދڽ(���/�������:v�{�;?d|��i	�Hwn�qY#j9�"��J�u�S1�0t�^�x��9|���K�+	��/��cHk�%ڈ�q�J�_
�����E=�TW�n��}��0����lEP�i���Zme(��S�߅:y��/���s������Wd0�h�Z�18����t�!Yjz��!_���[�����}��xB��s��*Ǉc��G�Ǟ<����f�?Be/�I�G9�ا��ă��н�W���}�|�#���qǎq�O��,_ZbO��
C #�BH���������%���0U9��\`s���~ӿ�h8ҙ�J�&v��?� j�6����Q$(�	�Eb���^��K�<��������L�����}�9D��i�M]����5J	�9lm��3�sb�nx��&����C�(n����<����L�6p�5�kg.����lߊڳ����#�1��5|�G�51�f�bЭ�#�>Jy��O^��F�wMO H��u����is~|��R�Ty'�����<�(
�ԃUUa�K�l�Υ6�,��R�(�@�ߝ��3��%T4W���e������n1D����!<�:\Y&ǻ76��ҳ���GTs���@E��2{�ݨO>�Hg�%Kof�����)�����lGJ屡M�z�r�t-�J̯��~)h�"¯8<u���+���̸���1��D�	��򱵡����-*��\���j���/S/�Y]9ɰ#�6}�Uo#úBSE���nn�:��+��V����K�+#rW1om'PU$V�b���m�"�(:R�'N��'���i��	���t_���W�;�����>l������g�q����|��]�٣oϝf:�t�.<��o=ŋ��K�N�p���g�[����{v�vm��?�3�|�5��i�:�(r�J ����@>yhޣ=Hߔ��J�C��5n V��,��>XL4Q��h6�x���O$��%�4�(u@T
��#���H�Z9��ӽ�:b�E%#B+���R�D$I�T���9{�ǎ%�2�x�Evڇ���c0*��J���,N|������^��8������4zv7�o�qz���2�
�kgf9��'��f�SSa���V�� �y��<*3D#�.��	)����w���?ȩS�������Y��i�$A�I#>2�����Sy��1!�I샢(ȋ!�t�Q]�C�K)PR"�d�`�B���}�vBnFW��_�������W4O%�5��ʟ ��a��O��.�$���r<"�E\�-���'�F#уj����-�C|�[�r�4�Jr��_d�C<�[���$�����Z����Uh�VA�zD _���ß�� ⠮��2N�� ����)q%����/>�$W�0���K�����e�.��X��q��#���wh��:b�4 o�ҝ�J��#/+ƣ�Fd����+�|���tw,0<}��;�ZK�2�0�R9YCթEL^%���}�ʜ�L��x�S�Y~�Y���>̾B����������L��;���'X���dS���>�^}�7��^���P��]}�5����5�����nv}�	Z;��ܟ|�/�F�J�vz��&�i�'�5�zr	��)b���D\n��E���ؼl'u�v�O�eB�C"��3
���� ��V�h�C�x�Zc�"d=��No�����,����ԞV����w�@p�&6��S2��W1�m�����L��I�MD�4E��G2)���4J&�v �R�.����#��� ��w�~�Jx
	�W��O>����#�lE+(� *�
�G@��iK�Mڴ����d��6֞���%��`�dCS�驽�KE��W[\��G��Ș_Z���.R���2�ᰙ'B�i����L(���cb����V�	��×�(tosL ��?�c���-%�p! dDi���H��FcC���<KX ��1�c֓��]�:�&��(�O,Տ�{�U�U��H� ٞmȱf��8�gE���0!x��:�XէPZ���E�%��K��b]d�ms��ˊ+	��F�ؖԮ&z:up�{�߲ ���cX��Z���Z�5�XլU��]W���Mt�����}`m��N��2��}�s������gf�[�sN������-��i�۠���LH�w�f�|E�2�3�L��_��^e�ٗ�����m7�봹��{9*'�x�+��Kop˧>ŶۮE����w��ŷ��ۯc��7���~�z�G|�����-�涳㾻���6�޳��_f�[����3sD��:��*Ch���S\ψ)RҎ�Ư%!�fMU�'-�H�ȵ&�\�j̰��D��\�·Z���L�$KE#�(8�<�!;p Z9�{d��JO��҃&-xqCr4UZ�#���?�o�k��8p�x�a�m��?w����D�0�	d^@�M���}����a����_}��C�@E�ג�S�;� QF��tAR2	!IĨ�v�|#���<c1Ր����C�yKiK�n�����F���P��t�]2cWcʪj@x&�օ����Ȕޠ��k&3I��=s������ }��9J� k-J
�fl`�B�� ��D�`��Iu��F����l�
��s�P��*z�^����α����C8{���i��:�]Y%[�"��� � L�xYz���*
�-��l�W=�����ޕ*�W�/!���g	�b]��^�oY��2ƭF�����c��;��x����Cj!����q�L1PB)��9�v���Y�p��gk�NA9X#G ����m��6�-��xf	�VPL�.��Ji��ee������T�3_tY�a���|��'�7��=��_r䖛��5\z�4�~�Y.������'��շ߈��g�0�kw������@d9�l߇޲��`Hw�~\����A5X�S�������^~�կ��'���m��C�j� D�Dђ����i̝~�$���VR��qo�"�L���1�R���o-��Q���h����-[!�Tx]��S��}��$�XH�u��1��B5z�����|���̏�P��{���' �r��kƾ�e�O�
�/�sT��-��d����KϞ�س?���nEd�"3�Z6�(M��h��&5�e-4�Y���o`��w����v
����|����V(�6
OpdL�3B��t���kk����"������e�&�����l��Z��?7BH��R���Ae� ��=���Q�(m��d�+�x�Yc�[Vbͮ�����cf�N��3��#�^x������s��2s���u�X�_�
����##�h)�K���?��G}��Ħ������}
A����-ڻ����葷/x������2}� �/�:Й����#,�އɻ�uD�-\�(e0� +rd�Q��`�"V�u��h̚��^��������~����y
[�E�rMdy/�(:���FK�Ժ����2g=�Rr�����o�����'�s�u��n^}�eΞ:�̞m���"�*�=;0[�F��t���󟣎�-�����=����6+�>�C_|���D��������˿���g����0�1��,���(7����l3�����$t!R`���kF��jK��Lk�(�)A1�Rr��p.9[I-��+n~�!�C;'fiYTh@�M�M)��:���"��E���Bh��`4(��Ј��QHs� N$�T�B+g,�]��=ݢE��\x�-��2zf��Rg�,f�k��mf�&@��D#����f��s��W9w���B	I�(�%^8>͙9b�a��ȥ�nbdT����R�x���
ZYN&*6(�w)����>�PZ'�`H�� ��|�?�s"�D@����!�$���"�<#k������X���D���2C���h����K'_<M����tۈ�cg�m_p�GzZ~C��1R��c�gZ_I/��"���^�	!P�x�I_�屏o��KIr#�1WB��ŉ�eZSS�ڵ�{�u�e�Ϡ�.E$#��"�c�yw�Q�`�`P՜^]��g�^��-���C�E �1"�	AЂ2��\��9-�����������"�x�,�p���غ��k��y�_��8�'E<~��ﺕO}�	�w�T�liT����q�{�`WkD(p�?���������-~���玞�?�������}V/��]{��������䘄�V�ˊd�D�IT$�o�hDSŅ��FN J�ih���QUQ�պr�R)�J�Ab�A	Ͱ��3�ĩ�G|�A�|�A�@I�Ҹ���,hט(��H����Q�ƤE�[��A��YʺƓ@d�&	IN��(A��`�@�R2���'�Y9}B�+!���j>�:m*�D� QJB��C���5_�<����P�Z��`T%*�-:6��J�.Zt�:����r.}~eJ�������B��\E.m&�3����9��N���,�ZB]������C��u�Udxt�u��#��f������y���|�+�d�� �����a�<��P��t[��V�Y!������$��a��ꟻ�ޏ� ]��ĕ��8g��������:�ۼ�j�����v�`^'����m��C����g]H�G�P�Aꂢ3�sP�-��8���fq�������݅+.Wx�Z�I�+RiA����1E�<���t%��K�wNS�����ұ�hn��a��yN��?������?�4&xTb�P��\�������ʏ���(�	F��CV{�V��-�p��p�=�s��Y������_x�ŗX۽���E�W����;8a��"N�P�@�HSAOZ�0H��sLT�&�l!�$^�q��'G�<":�iOO15=�L�G���+r���bm�;wp����ر ���T��F��$��$�My1Q�Ԅ6݇�i )׵��v���iF�?�2DT%�?JȻm��x���sq4��#��2�_{�67�L��D#Բε4�@��U[9�Ç�r�M,ͨȩLF$BJ����)���E�V^�e9Jg8)뚲�!��������t�ul�F'���~b�(�8H������&��w͜���IFXG& ���J\��$zǅ��8s�,n�5��{�g����s�t�C&aF�b�`�~ G@E�Fϔ6�!�q�'����𞺮�!*��˕{t{&�NU!�@���I���@DJ[�u�D�v�,GJ�ݴ��q�b���"�e��!|�,*�<���2�w죘�f�ri-m��k��:
Њ(eFI���_q*���=ByT��Uɶ"�J"^}�s�?��믲����>��=�n|�m����|���7�<������XS�#:˸p�?y�yv^57�v;ϟx�o|�i:�q����o����s�ku��'�!����zg=q��D}c����6�RJ0�*F��p�sZg�B!�D��C��m#y��%i�{=}�1�n���A�\�>Χ�x}��^#ʈ�2Q�.To�<����.O3�G����>&��L�z�DM���(�F`BRHM+��y�ٗ^f�ٳLM��D���sD[!2IP`�GɌd���SpYAt�|n�]=�K�O���Gٚib�c�T^����=E�e���&ou0&c�|���P&��{�9"%s� Ҵ���|��Cڨ�������2���c��'���'���R��<�yUJ��j����h Ȁj���Ɇj3Bn��1�E$
��0��O��%�O>����`v��j̞�L�?���3�(�FvB]/0d{VE�BWħE��C��+)�W��/(��ܣh�8���(f���o���qI$�2|9�*K��ԃ!��2v4@��(S@��6��<i��+��_#�e�����
�Q�Lb$7�1&+0E�s��5K�s�Z9Rk�AEm@L��D�_[�����h��kG������C:�ì�v�$�ϝ��7_cǃw��������/�=7=�:'^?�S
�2@��%-�nN�q�!o=����;\��CZ\���Evo�y��پ=���[q����9�#��}�{ O��IL��1ѿ"`�Ë$�[xA����1�Z��,fi�6R,�;�ܞ�z�Q��4e��|gM��l��Dr��%Ȑf�"�;y4�f��+46��N���6��t_D2�Q�6��'���6���{�lՒi���!.�0�����S����AI�Q
Q. �l�{�zH$��$Q�^hL�f��av�q'�?����b�G-r�#�����ֲ�c'FgI�gf�vߘ���QRbbR����;1!�����h����Y&#�6:H1�'H���pv{.'��Xw	l6]�8��������0K�,��
'��;���Yf�cFD��ef;�l���y�̙L?�r�àOCe��x�r��+��_D\I迠��1X\=F:���w.�������)s"
EdFF��S��F�s��[h�����&�[�8�p� �A�D?��>���Y*��Ӕ	@���0y���*2�kfw�?����y�A����m�s`v��%�$U����BM�#^�nL7��Q
�嗎r����ڷ9��G���f���#�
�Dʊ���q��ٺc;a��9��|����@tZ�N_�������?���1Ӈ�3�����딗iY��V�w%�w-�4��bR銁H�)���`��&2v5CW3�
L;C��
�4��᪇�>��tA��3�A�{�*ـ� צBr�����\t5E�j@h���S�MU�h@DD�hrD�hd$�M���m�E.[�:����1}������@z�β�����iL��ВPG)�K 
/23;ϾG?���ĩ��!yn�bzD�	�uI��'zaV�%�j15=�x<D
A��<&k�j>L��9��_D\V��͝�Q��ύ�kN���ݑ����������p�����׎��s��.2�m�f
���É��'��SNr��[���y��+#o�((��P��{�<}��QǕ���o�Q��[��E���o���9/Z�آ�*��2���/3|�U��e��fi�˧�M��=���G�_��ה���"�#��B��#5:DL�b�6f0�	�E{�N��G����N�%��U

�	>2ۙB�,q�	uM,Q+��B�궓L�������:�N��<�,�������'�������:�V����[��⦽�����_�Ƌ/�Rm�~����>|Y�U�N�Bᅢ%S�f��2�ƷHT�7���U>6��w/���1&�t9_��4Qz��/.sh�N��`Z-V��w�;﹓�*�Y��*U擗���d���Hl�꺮�z^O�%g3�:.`㽫�_�'����EH�*m2$4:)4+K��d�0`��I���kKkt�WQ�CJEh��ξs�?�w����2����)��v;��N�J	C!Q" Y@���&�d�w���>Ο>�s@W��
���Q2��[��y���j ���i"�D+����2��ːa�n���m�RE�8v�ߙƸ��7l?;�,�����ǌ��$��k,"�.X��̎�n���Q32A�,�O����b��4��ـ<�����*P�+��_P\9ʿ����{ʺ�|&���_��MnF)r���"�^��S'�~�s�>ǖ�).�������B�
��-l�=5�s��K,_Bǥ�g�$���W8ᑍK�afj�jXsqq��3ͭ��9�$���?a�[B&ie-����1F	Z�iZ��&I�r<��F��PA���EM��K�9����aO_r��y]�{�W�2s�ut�6�S���K��ԏx�7��S���g�㈚i�	����@�(<��d[�d]33oVl���Ш�5T�w/�RH��I�;�*}��Hf$�n�9aYY�ӝ�E��b�2Cj�6�|�ĝۨ�@L�7�ԓ�Y'�s�&������"��E����߈�"7��ވ��7Ӏ�l�UEU��Bc�%GMmnmD���gO���ST�bmq	_W�6QDB�D�A�v�Py�2��{���Z�^y�� 	R��BH��I�6
�p��l4�OK��^�h���D>��.���!bVL��ɦO"�H{ӟ�}n`�717�SދdW��'J⽣g4��U���t6�jϰ��(n�I_����	.��u�0[g,��!2-�̐��N��
B��������������=��<BW��+	�#��>�Ā�K��BE�e���W;�ʖ�5�,CuV��*�f�.����ѽ� �{���_^���W�CD��S�ߠU���P�#�� ��.��<'KP�+|�*��+4K��*�Vx���ا(���3�?ˉo~���sLIŬ��B���v�� ��,WC�L��tlы�ve����In�TQ�1e=�u��e޹x�����Ǹfj�z�8r�ﾋ��������Fj��*��5���x���F�mՌkB%�XS�E^��oBx�F�Zl��ߝ�'-N)q�L�k�
-:�hu�yd��%�����tn8B�k�1$��f���5Jpoq�w.&66�}Zr����m6�(?\���X�tT�~@G�>�K�!�J���*�y���؛o���9z�v�b�:7���,�r����R��!Y�E�$��
�O�����<����7���0���y��ߺ��s�.�]@jM�ߧ��R!D�0eJ�c3�;^��/��v9~ٱ����X��덝��'��?���z�gr$֯��WS�f̢b ,��de��h�����7�N�A���"�g���U��T2n�R]R�&AxD"N�1��W�[>��?�Ȕ"����C,��,���G�v+�kt�V�#P���ry�������G_����"s-E!�n����ڍ��_Y��+��Z�g�W������lv���C(�G#�ѐ�����Z!�|���#��ĵ_�;���#���o�-/��߰�Z1���t����9��`����vyI �UB�k������!�^���x��'��u;_�¯3w�]���a��wb�
���:��*�>`�J-uq����gp�*�I-LZݒ�,�z]d��*��E�B�UrC�U�qt0�0����ku闎se�j�n��z,l%FIFF�&	Ҥ��B��^7vZD���"~�M6�y�9�o��'.e�o�[�]6w?y���Iڅ!kZ���s��d�|��Ko������1� ;���7�/�W�&ƈQ:i���I��sҼ)��p����ݷ���������l��3�刺�����L���
���F c@�d��_7ع,�m�ԣx��-���a��R 4-v&�\�R��k�������˻*��#s��;�Vj�p�v��F�;�F�{?��׿�����ؿ�x��VF�,��kLO���bX�kMm���B=�C|Y ����>��~�;�p]��3�$�0����@L��T!�����l��Y/R�P(a0�-�+FQ�d�tY|����o��x5yO�u2!X������X�u`��քآ�.0JQ���P������(O�c��E����o������O0s��L�x-��n��?�Kμy���k�{�@�%�yNɥf�gA��ڵE!)�&��4�v>�0�* �ǖ���i�`�[[�W+��%ܝ�ӹ�f�LA�₦��5�:U,U;��c������<��K�0=���=d��AD��wyY�@`�P״�-�:]�WV1ZS���r�^۠����(�b��i�s����_C5�j�{��<XO,d:U�ɿ�PZBȊ,�V�����3Ț����D�`#T%щD���6��G@�	���������E2���!�����#d=�+��
f�f�0Ծ��BŜJ*�C�t9`��gXx�>"�Q�a��� =�$�w�j\���R��&@ )�9"�d����������SN2k�a��r*7���Uy��Q��U(BS�l��6��o�:�rl���i :�� tyč��~�'wX��O�AA
��x�8���Q�����41F�TM%../����7F��Կ�SE�K0��ﬢ��c�����ɓ�����G�n�b0�kkb@'q%37��y�e+�����u��_!Ņ�#>�uU�+��ĕ����l�����������6��,}@Ҵ@MN<�4�����r����/�љ�"2A�!�e�aY�Sd�R�$��`�H���}Ğ[�ua�^��J���C7�J)���̳�����,ӷ�'��΃���7��'��?�p/3v���-8!��q�w��R<cb��U����3��6�`T���u���θx�^���=�U?��b��k�y�4�&�π�9�5yt�ӧ��
jq�))Qα��'zp�#�7�h1�u�P��>R��]aX[]F���ͅ����g�����O��d��jZQ�u��e��fF��ړ�y��!!�F ��%x��k�F�u �@&�t�"4�.#B���d�F�tj���lrk��&�E �H.ي��.�sj�i��k��Z䲅�ZD�\�Ƽ��3Z��w��
�!ր��"A��!��/k����	��uǽ��y�}�;l����]:�FS'�2Ռ�dZbd�Y�\���?L�=�����f������6w��t��'�o�d����[I��E�ZHѢ��ŷ)�y�G�T9@�k�/���k
��@�+� ɧrD����3���>7��S���Z1"����^��}q%�D������ҡ���ډ�sU�g.���ThBIA�e��WV�2Q+V�,�r������-� s���=�r���"Ԟ�ldK�K<����%V�8Evn�L��FE��p�����=�Y^}�N����^K�}�j�۶��;n��O����|���"Ӆdf����/+��	�R�J�w5Q@Gg�Q��;M �z� :&gG�\:z�7N�'��,�}�]w�C�P�,�G2��O8u��_��z���1%:6���RN����}�d�R!	֣���CIY�ɕ��*� ���na�ݷ�ھ��=���q�"ɼȐ$]�M� k��!��ӧ��}��AhO��� �ďP��Ʉ��>I��dZ�uL��JT����Žn����/S%�����".X:~�9a�b�:U�:@����Z2�n�x�ay�{"l� d��(�]>�@M�DBD�$�S�o���<��os��Q����&�����h%�E����E�e�I��,}�?M��Æ@c�uc���LyK��WX|�-��"���޵���9t��t^}N�F�y���UzJ�Ku��i�H�D�d�C
E�]I;U\9�Q�R"���DW;񹕱�uW��r��ՄB�i-�CE'+j��TF�R�r�-��/���#lۿ�v֦��D �Bc&�Ej�w���Ϋo�^>�܊��]��X���R�QS�,�����Gԫ5�,m�2��w���MWq�C���8��숒���?W�#U�F��Y�0�&o�ǈ����K,�#����#�*�QS ��k����ko��̷�����"S�݉�y�amH��?��O~���7).^dNI
!���)��I�%M�Ӂ�T5���T�gR�
�f�]�)Rפ��f0��z�u��f��� �!�vb�	��cL�i"���9��7������~�#�<�,�|���~�Gو�
�h�]�Fw�.��YD��u�PR�7��$��ζ��ܤH�$R(�>���l��'��HĹ:mPD�@0�5��s���s�0B5K���f��BD�.i+Is|_9��	��-[o��#�=�;����Ӥsm -G�B*I��%:�e4���'�GN���_� ����Wx��A�6H�ʂr���l]�����UO|�b�n�v���o��g��g~L�?ff�4�]�_c��u�Ǻ���W�)b���R����+U�?x\I�A|���#bĖ����p�����t��uIK�us�͞�@��5J+zy�q]2*+��ҕ�N�3\s�/�x�����Aj-������b��"'�9�9f�Vљ�J���1��<��?�S���&N�8��{Rk��*QTa���{7�G���9���q~yL'j��5�2�;Jg8�c����(�aC�����v�����31ү<���8��ęg�K��1���:�z�M��%�MF�d�F�
&���Z�q����!�$fH�sJh��T(�Y_{:���i���-��e��;!��=����I���&��	!��(�hD���x�g^z�p�oF�ޕ5Ξz�3'�q��y�����c�`�;C��"{�^����c��kP���r���>���*�\`�;�u6�i����(h���Y�h����c@D�RA�'%;�6'�{>�iD��.�
�*m�i�(�1���IjV�4���S�@f
����'Y~��>�4!��9�RK�b�9^4�"D��<wx?����BlJ�q似ɷ����~�H�H���h%�H�1��#���V����A�s�Os���i�.1X��ҥS8?ffa�p�"�P�s6\���*�U�+.���+���&�$����'E�HpI�U�8'}�Gy����\(o��k�!�I�9ޡ��B�C����#Ɩ��4��93mB�PqM�3DR�V�K�d�s7_�`X��s�q��r��Üz��y�^�ß|���߆l+��>:DB������_�9�v�����W���9p��)�y�izs��i�rL�jZ��;��F�H�ɚ�r��&j�ؖd��PB�
D�(e*�ЖtQ�t�(����u�F����֝��ib=�Ā���B]>�l�O}��IC;�@�l8��@n4�Y��X�V�Ee�vÍ,��O�f~2�6T1b}��,�q�}"R�xHG�U�3��+̜���?��p�]Z�P���CZ���r�>�r��N��-^�����>q/�O>L{�v�1�2�(Giq��'�o���?{�d[v�w����>�\�73_�|��+o�2@U�
_0H�)Q�ZRK������111��L�L�L���F�բ($R  �[�T��wϛ|�9f��}��|e Tr�[�2��瞻Ϲ{�o}Bi�ٶ�_�5��GI`,�t�1���u͐C�!/^܀��a�"�Sg�����1�򿉉��K6�B�!�D����=��?�>�,��-��!EY��X[0���<H����?c��2�����)��1I@G"���*6z$:�Ƒ/-Q�t-uϱ��M�z��jT��t��ǘU���1��)�V�0{V�_����E�l��
�7�����q������������ly��@�2������+���d�	;�d��q�.�.Ê$��&�l"HL�O!*���z9���z�"3АT�T��a
�ِ�w�毰�{��>á�������#�X������#�����.X��	������/|���}֟{���Q��_�,��G��~�������|��_�g�y7k8h�8�����Dm0��L�g�;�����\
qd�"a���SP�%�XL��'�4'BljL�Je�T���P�뚘9jj�L\
��py�XdLq|�ml��������r�{>�?���9�r��EȜ!9�]����^��j���nd�+Y�7��-$z��Y5C�g8��� �*��\���'x��g9��ɞ���`eꚲ��u>@�SGd�K��\Q�.[PiHr�
�����K�Q)D� �1�to!MH��@��4��:9�`L��<0�Cv;�n!h�� 6���P�j�^�45W�w[O��ٿ�2F
�nq�ID	3����o�I[B�����"	�ڍ�a_���m��r��4?o��A��P'�M��O<Ovx?~k��ߎ���E&�1a��g�,,�pf.g��\�.�5����A=ރ���{����2��O�.;���}�c����i�E�?oD�-��1mH&����zJ�{�����!e��s�5b��P�HSz�(��M���B�0���/N`����w��,^w5�c��ư��M7��X�d��x�_���O��������U,����Bf�ލo�ʃ�]y/~�+��o��\���7%Lkz�� V1���I�'�w��ȈM���$G#-mi*�Z�|c�E{+wf����S{��q�}�ðk�;YU�Q�T�*T���v�bŉ�-�m@�K��5�\����o��i�0������ŋ\�4�o2�j��l/�CU�
(<1���SE���0�ʩ?��_�KV� ����3�j���F��8t���+X:vw�,�`5b�>{8{��?�J5�D�3	����#� ��P�k��(Ӌ�duCh�	�����
�T��8�ͮ�k��l�./(�:X^�{�ɣ�}���-V��X���{�o{��]���%�b�-��z���ZK�����2Н�Q'�B 7&��-1ǥ�_��Rb����\;��_�%�������3[L֞bT������.�.��꘾�Q0�1�bc\�gԓ{��gU��c�h`�UA�e���e��S�Q+a�Fr�ᾉ���_��рe��q�y��,�+)/1+g�1H�o��c5�}-vzh$��`���6/���ȆK����x-�z�&ۻ���W�@��8���x��b��	n�孬4�=�$W�w��!��!���_@�e��{Y��&��f��/�Ǟy�c�>KYNӔ,�g��!���Y�]�%T�툗1b4iu��PS�ow�P��-pH[�W��_�Ὴ5Lv����L���Ǯ!��v���7��?�������JjH��&��O�������H}�O}�L^~�+p�~J5�b'��	4� ���qL�`�a1�Q�����K�^β�!X�B(O�d�GЅ�+��x�u�q'��W�BUS�8N>��x��vi��54���GL� �r�&�^��!9�$�jZ``��匶\ZEN:�#���+������)�A7�Ѡ8ۂ_��.ۛ��@�@����*2~�	�ߠ��;��m�~��X29}�ka��J������iC�0�?����Fl�5j>�<�bNZ��=�Y>�����/~�?�������d���n�8�d����G���z�猍U���7ȎW<�B;{���J�U_2"dЈS%��6_�"5��beyl����'�{�C� ������s�}� �9&O=�ß�C�=�C��"+{��ٿ��f���W#�Qp��������I�h�{��o���ȡ�~���;��o�g��uΜ<ξl�(TloO9�0`����1.+�`;'M鐼��`����&!�S^H�=�$'w�I���+�>'vqE�wT  lO���Y�+������[��q�M�C2,L*����tھml%=�v
[c^��7x��_�ڠ��C�3?��⠗d�$~�9�Z�#ۨ�ʚ�I3�2'N g�5���Tư�q���l?���'��C஻�p�'>�Y��IV3K��Ŀ���ZS[�8���o��1��YbPPA�IB,mF.q���]�C��[�@MDQc�k%�s�ѻ���r��[d�����r��|^m�������&e$�����.8"{l�l����ט~�a&lnM�.s�G>ĵw߅�+^���g��y�ڂ<�)�F��M��3a��E	�2��֪�j�S��T��J��l!�0�B��H/k�=5����fc�
L�������/��뮥�iYw���~�$k�u����Of���Y�DF����Ӝ=~��G����\{%W������������:*X?��>�}��1��!2�KBb(+Ϲsgy�q�-oe����4���p#��|3����?�ǜ|�A��5�T�=����2RW�9C���f>G�.��#-�&����.�́�,��G�?�t��~�����2ǃҿ�V�z��HYFK������Er�: M�#U��/�z<��o���9�B�)v�1Y�@f�!��-�zmN�T�1A�:uKe�g �@l�e�D_B�P������2{�	Μ?�f�]�Q�moaăied[��D�F�Fħω'��;zWM�v0i�]عh�$�";��b�.ȅ 	LWFC6\������>^��s,, nV��q�=�4����xk+^6�UFQI�Ig�a����t����򞷳���#��f�u0�2��&.����bo�"���2�f��Ս��t�cQ���D�����/�+��W�?{���
�o>����T�&3���P̑���Vq�X�,�������1;N�]N&���y�K�D�kk�o�r�,T3�
Y���Pnnq�K_��G��{���>H�g���q3+�et� �yl�a�q�Ͼ��b��UT��Y�--rh�����M�������x���_�U��{|��<���������>���j�ҙ�;'=Ml��]�����ҺAhEY:64EZlw����U֭S���2�7����\���b�\A\��l\lG�2K������n+���)4�����&/�b5/�cC*�~�4�X;�5�7`�&q�Gݹ�F�V�}���X�;0JK�@o���G���'��&�M��D��듩��B�
�@�ڭ]�m�n��N��Hl���K�'�;x�p]T�`�b�e��8�����w�N���~�	�����/#Ix'�֙M_��N�M�I�iDCJHBB>*y������+���v����%�K��Ǖ�y���}�����z?u�Ņ��b��]��v"OB��5��˽���]v�?�Y����3��7��Wι�&Fk�|yf��U]ݑ�϶����n�t��q��>�R�c�������2�(��B,y������|���)�ﻇ���d�[�K��zw����s�Ĕ����L�6���ٔ�x�J4�����>�g��y���S�=vq�u�(W�x�|������������@�ȣ��#݂�>�i�CM�
QQT-ARy]�`:g�-k���F���[31�ERf�\�kE*B%��<��`���f�<UM�`2���i<E���2M'(�(mGZAC`�ŗ8�8�(�^f��M� �1i�!w�K\�k�`=5��&��>���8��ǆHBB���`�
�{$z��V�m�$��L&	�fv���ɭ�fj�$u7��Ƚ��yt���.�������s��u�ܼcx�����SO?G�5�@GMj�H4�
�)���S�u���Z�[>�|�^��_ޠ����>̜���i�ֱ{��MY0�o��]�=T$f�l,��Q���� ���~�'��8�n����w�����S� 1���)KK̪�[,O���B��H|�Ơ���\�O�.;���}��>�Q�ijrU1����זL�2�\�1�'	OHWߵ��f���(��+ە�i���=��v��a�7�$�oAP�)ĐQa��G��ƹg���Y��~F�ߋ,�{�>����� ����y��}��1�<����i���C,��o��Qa��1/=�8��6������š�n���ţ_�,�b����{8���d�ZB4�h�A� i~_��� �f�;��-��,��B깶bj�I�)��t��^Q�����7p�?HXXh{���<ֹ$ߩC���;�N&E�"�5X��^��Pk���D��dPm���'c2�al�^� !��i��
Y��>i�+�L6�3�{���"j�Ĕ�k���1��V�6O'��GZ�Ym@}H����,UPb]��:۪�Q��m�����6Cw.�n/$�����+���ӏ=�K��KF=��U�U��D���Cb��`R`��'b�,~Lm5	mn]
p�a���c粖q���ҡ�_�^�q��!D5�5�3Aj4��{E�꒘��r"�{k�M�1� �+�� :_��?������-�bBً�X18���6�w�˅�Oqq�qJ,��G�ED%�	���4B,v\�����x��pv�=֘D����	��}�>��_xC�}�.����hN|�4�	��C�w˩͂��!�#jĸ.�~e&�����.���gN+�� ��]f���Ɔ��NiE5� ��ҫ��~�<�}�Q���i�|���cL�ѷ���w1:��_�T�z�eFα��K���f�U�ۮ��<w<���'��=�^q%W_uű��}�{Y��f���?��Ğa!��l�qM���	s`�I@(<�4D�1A�a'�ڭ�!����:������d�����`L�1�`<������
��3^Ye�`���h���5Ԝ����SF�:�-C��*i1[�V�ct�0���@��&6������S�"412mRE�oκ60I�m�1��4e��G�`$�"bd'84����J0~:� 9��J�k�}WO�zg,݇*b�����zJʖ;V�@�	�n��i{ݗ޽)h����6�4� }�}G9�������9ð�&��ba��1o�hQ�S+���$jGtS�Ƙv��2mj\�#�!eM��^�Tv�����̐�HJ�J�G�0"�:�D���O���L�a��>��w!�w��L~3h;��޻����xMM^G�Ʉ�Ԅ�՛����������O�u��{���T#����Flm�ho�4�o��}Έy�4u�Xǧ?�A~�s��N����C�+ا?�a$��dAm�M������M�n[��e������.M�y��fן_c#I�Cy�c�K����I+\��='�L>����s'�?�a�W^A�_P���L��1`Ze������ig��s�U���7�˧>�/Y,q���$[ڃ/KB?#��(��ί�}�a�~��YE2a �+&�#6ǅV�O0o=�Hd���	�&�Z*�	`"E�(|�X1&�|�s�Qy"+�Y������c����1@��I%m�Qb ��.�VH �e�ګ����~�q֛��3��>d%>��Q���cE�	Y�aԶD-I���ib�%�K�ڌ-%�:�	��=�k�g�NtW��5�5q���XO%�QۭGW���$�X���4F��ړ���z'�cOr��`HV���DTЍY팰��t�$��# �,k/2����:��4](U�̥�C�)���Zѝ �ủ�p�M�)K�`���6S7���?�s|���9)����BV~����x;�w���'9������Y:|��6�̈́�+�(�DF=f��\�ίߺ���e��l ����\z���e��&�w�)�"y`M��sS��[!j�1��Ω�Z�e?�vm�?�^_�yG�������g�����y���q�٧�p���I��w����QB1dH���ޕ�p���(︎�_������|��=�<�����!G�x;Ma��33�g,^{%���_�K�=ƙ�	W��Ծ��˨}h���X�� ݜ��
�[�;>e�7H"dQ��S���FI��	�����x�,�ػ��w݃]YJ�0��u�T��&s���_�;i������t��~�v3���ٿ��F��K�Y��鬦�*bPj�)��~�'�PULl3*�9��S��Kh��|a�`dxٶs樲�I�%�3%�(8%-IL3�ږ��b#o��{R��ѷ��h���qO<�0N���^���:�)vX�������0D�qm	[�#���:���������<Gc*1�>/i�Ov�ho�% ���,U̪�B�K�fZ_R �8� )hj��yF������m�-�d&�\��_�/7i����~�����λ9���Q�Pn�ۻL�s��G���:��w�h}{��#�W��3$V��8˧?�!~鳟���a~��C�6�3$z���Yχ;�:|d%˖��4�FP���jK�j���'�s�d���;s�TuW%N�sж�i�-˨"qF"W�i9�������<���Y������w$��>@���ۯĻ)��7�f�1���c��(���op���ʠ���(ͤbAw�u�+�����Lmj�#*������#-i� �}�v��g��©k*yIi���jHLt6�v��Y�7|�����$s��4&�6���n��5�'��Uuٹ��2��[n"����锾1���l@.J?��=TM�F�EC�N5�QX����8mߺ}��e���rI�3?�WT���N;���a�d"�/Jc����X��0/��IǛ�$E��u߄$���ob���y�ΰ����1ơ�n	�v��:ƿ�T!b%�v�B/�Q��4g��L&Xc�$Fb^US�e�:���f܊�� �l:cR�C�AR[�(i�0�YGfm
� bb�K�Нj�%������U�k�h�F(����GX��3h���}��������x�SgX[�[�7bk�,5�F�c���&F$D�e�7m���4��������׆�@.��C8;�%֤�a���m��m��U�56�]�;�Ɵ�^Yn��-��Ec���M_%2��z�f��`�1��_|��}s�Kx�p�1���^�;�.<�"�=��u��C��w�&��'�u�2����1j�:�������g����S�j����i1D�a�pi�s�w}�ݛRٹy�P@�[�ضem�s�5\���� +i�:&Ǚ|T;���.D�*L��R�1�ģ(1z��y;7���<��Oq`�Ġ���g�e�=�f�oP>�/�����D!C{�t�ǔձ�z&3��O��x2��߅���CZ쬫�b��[�Aj��6�l��!���k{pi��&,��ͲĎ(�X��h���߃{�!�=�<��K��N-�=@̴��e����i|�C�b�^�3gYS��&x�b��,mwQ��.*mjo���l��MS��1��[� h� !0(z����Zh�mU�vNg�=~�6���X�-�#ɱ��S���m��`�}���u+�{d�C+�������1,��CS86��؛-/nLg.��W��o��f§?�~�������~��C��FZט��ۂ��c�VB$�%Y?��v���.T�1�u�]���ꮇ~�D��絾��},���T����^=�W58Qʼ��g�����0z��,�}d�\��5}q���\w3W��~�\}:�dq^0��1�FA\�����Kn@f=����G���Æ4��XK0P�@/�����;v=:ߍ��]Ꟛ��h�m����b��{VY��]��&�dm��2l[X+��@q]�swG���k�"F�ַj������_`���y�񧨧Y���O���Db�4(����rrkڤ�#Б֡&Pal牐(��Nw�sJ
l$���a�3��窴�>5��A��֠�&9T�4c�+K�,ߌu̇�3H �}ꦦw�*�����阬j�aT�����_7�scȋ^r������l6c8RV%�.K����^Ѫz؀���E��#uUcDX.0+K�r�aD�U�r-kTb�h��O]�]z�no��~���agj �(�����k�������m,~6�	H5��K/�C�k,/��u��ZiCn�����3N8-Q��e{�v١�	�"تI��W54�^nZ6��rJfM�-�u����J+��e�0�O�����q��ruN�5��	c t\�)�����,��8��s��jM/7���H�gz�EΜ>Ņ���G�O��[Y��(�_��`�-"���f�1�&�T�%��ϳ��ņ~ѣ�7�M��Ål�Н5��!�v��֒	s��*���ā��guQ�����Ho{�(W}����˚�ȱ�I�)*��3�,A��I�T��b��DMe�i]�r�[����k��?��W��(*�*E�`ayal�O �G�0m���"#���-'�*���$d���s�6	�ʑ�ʊ��C��4�J�2�nSP,�e����C�E���l��ێ��-b�n�U�H�N��9�%���ˉ�p�λO������B�`P��4]9L��WUb;;/����a]�Jע�y�x<��k����g,�K�iJ�!�Q�rz�n�%��lʬ��b;Jg�!���}��4MC=-��T�릥N�v���7�1�}.f|�:���W_�]��*�V�P�J���&�
q���g�{�.�xN~��<�����{履+{�]dOnp�1n��W1}�F͞�p�D]��rn�k���Q��4�<��#|�O/g�o�.;�7h����ƈ�=E$��p�vUt�����6�k���%�E��ߙ#}m)D��g
�w�_fg`�u�֠-o��vUk[:{��I2oI@4M���l$�H��{�t��c�p|��#q�}�w�Ȩ�OeҜ��C4�iSkf���/!�O��PQ�&��58���b��Ѥ;t���ՕDu�#���U1#ڈ�'M:F�LC�F��n{�;ɯ��2z�C��E���$��#�s�&r����h����^rNF,b
����������%�.���H�D6ַXZ^bqy���#�p���:���9bP�Y.`��Pc��ѧ6��1�����W�cqX������*�ރ8�&�<��F�!��~�ĩY�t�̡�����͗�s��lqW�[���"�eq�>��nN>�_x��VzH��Մ�W��3��3�N!�c�`��9��k�!�$k�%�oS�9��0&q$��4R�5�o6%����~�#3_{���{ߪ�)V�sXk���U!Iթ�I�K�ۻݲ|�H�V��V�>g�6`���}T%��#
�{��'^`�%z��́׸�����J��s�ޢ߳��Romᖖ�x��a_N��2�?�T��a���`��[��v١�Q�F�Ӛa��}�	�0���3��5	0"1=W5��!;=(�R��-~�����FVܮ����A�t���L����]Y�n����%�Bb!׀i*
"E�3�5'�3>�SO�`p�-���po�uIJ4ɜD��	�I��'�/���X�p[yBSR7S�Y X����c�������wW>wVlgc��c"��1�&FO�5����Z��xl:���J���>X]Nk����۱0�vDRo��sߨ��0ɮ�CAG�k��������}_}5���&_z��UI�����UL1�	�^�mm�ᱍ����E�j�349V���bHcv�l��7_�9�]�?����H&1�ՙe�˹�a�8�w���;�D#�f�g�]��W�_���.�n�>��␅�[�J���8�e���~P"���6�.�7�^�5����FŇ�3��I �,��1Ш�12k����#��&Hķ�!�4�`�Z�E�<���.K|]�! "ə�9�<O&$�`w�]�#-�M������N�������B�Ƕon��ybCH���9e�`@8�M��=u��������=W�^���t{�ړϑM*]E��UŞ�+Nl��sК�e�ӅDߔ&���?�~�r���e����?�1	��)��κ
�f��h��)�̒Y;$tm0-:T�Q���;xW�޽Y��2Z��������:tE	1��"�i�e�i����`�#*H ��筒��m �B�qY`�r2��dL��s�/���O���;�{����H�Kg�k���l>�?�������ڌ�釀�T��i�wx*Q�H4m�^sGޞq�(���P�Ė�x<����#yκ�\����⮹�&�X�eMn3DF�e�)'2}�ߪh��f��B���4�O� yo:�ɮ���V?��w����E�Ν楇e����#TES�������.\`��:W� 5@ʿ��8�M�'J���IN�:P�����qs�u� ��z4�Qz�1�3�ta���(W�v+�w�����#NrL4)P�nC�j�o���;�^zЪ��v�r��޻����?���O�(�B��;�0$��|뜫�[��T3��#D���� �kFE*��lN�cT�T�.b0�$���ą2������{�錪������作�(ȳ Z?nvg�O�������='����#�cL۩s,@f-J�L�b�ϝ���u�CI~�lh��w����n����o|��/��<۠�9%?��?�2+�E.X�BB��\�[AX�
�i�{�[��v١���/��"�4"�RV�����e�zJ>��1`��є��^�!�3����)ki�����c�H��D�m)��^�+,�DS��h8�����ї��j���E�v��zIऺ-/���H$ǐ�A���f뇏��Oq�k�`宷�z���!�����y�_%;~��&�EY�5VR_3����4Jg	�y�Tf�4~icbg-�#�-4˶$f3	)��qbs±�?��?�1B���ÏK�<�8��2���Z���l��_�F}wɄ�n�Fӭ`���,��3��{��������a�]�,�Y�y�F�	1�Գ	��S��N�O+&��p���(Ϯ1h�j�G N���\��4#v��x�DJ0B,zl���4}�{�3��
��z��L~�����Uq1�TW��C�i<�MX�����-�N-���k��n{��y7����l��@$-r�R�A#�L;� ��5�? �w���t��kd2�2�J�3H��!abl�W�b����nF���m�]�`��Y�`0���C`6�Q�%��1X��E��sk,�+n�]{@�� �.M~t��w�4��Vg���D���'�<�V5�e6��l�������=@}���#��87�b���'>3��җq����+,�s���3[�,.��#_����JL���������nv١���[�&��"ƾ	�*k�y�r6.b��:�z�6C���M�עŰ\2����s������[2l��˺����)��+-e��k4b%���/cl��wN2E�O�;�:H�� &��ՙ �A"�B�d���d�MΉ�=��Ǟ`�O��hq��p�/�GO��ڳ�(u�L�b�oRV^8yF��4��i�J����]�k��U�ޝ��1j�u�Y����?r�;>�1z�0�<C���A����!��CH�]L�՞�������:�Idf0H�@.�6�Il���C���J�� &�Z�A���D�5נwO0"���=s���lN�x�E�?�0v<e�xdV���:r7~�(j�1Bca[�����+X�w���},_u5�ؕ���4�V�O�r��d�zfCZ��f�vg�hd��}��,�7(8��{���wh���!h"z�1�[Kٔx"�A#�5��>Y��X����E�~�p�"eYb$	+)m�������+���Aǝc(��a�G�1����U�ϖP�ZK�+p.K�QL�*k:JZ���/u�:���_z}���_�����]�!Y���R�/��������V(�<��=1�s�~�ny����w��3[1�mn@Y��&���Ui�9�5P�%�?�����?�܏�y���e���'�c) n�b��2���8��|t�>�C[PΪ$x�r�Is�����m?�끓���53��)G FO�Bl�-�)�n�ҹ�
���n�y"Tu�AȜ#s�uX�L�����T��K@��+�X�mH�Զpڕ��1��%�A��5�B��~�~Q��NR��<�p�ȸ:/Ȳ>���̀&B�gSO3*y�f[�$���Ѥ%BL�ˎ�)H���=�iKA,D	ԍ�܀<_`b����w0��&�rO�EF�5����ڔ5I�ׁ�i0��d��:5��K�vʘ"���| ��r,�C�=�<#�V]΂YZH�BU��"��A�����,'3��q+Ҏ\EV��_��-�ŋ\<q����Re&xLL��8��q���{a��k`e5��q�롡I����F!G���9al��c��^�:��h�R�&�=@Z�jZA���7����/�'z�oP��-f,����m&���éP��'��WlM�lll��9G��a@�Y�Um '-����	a�}����U�{=��>��x�P�%�Y�zqi�܊�pE��[�C�U��x�9�S�%:!��&���Hl�����& Z�Y5ġ&e�Θ�5�s#ņ�
��=�}Ԥ�Ԡ�cQ���ĳ')V�؅����iο��O��*�z�6I{�7���g���������{��i�VZ�P�X(r.ۏ���'��ZL�ؠ��HB�`&���rRh����x��Иf�%ω���b��ݥ��� �o����DI���fBM�̰��4��&mz^#>��l�C�J#*�!�d��Qq�#uC.�,B��8z}��X�
�
.mi�qyK�4"1�>'B�n����k�Q��B��x�In� �^ɳ��D�����`�7$�s5�8����J*v�-�%|@L������&�3Z�� ��D� ��@�3�l��%i#�VSv҄�~ev��pmScB��@H�<I����뼲 .�uQ�cmZ�L�J(�˱^���IH�`�v��6_�
>	�ā��2r �V��c"���ե-��n���,�1���<�u�$m�E��]M���q-�.����6O�k��;"�:��@�lrjѱt��y��_���f9��o�z��P��ܦ�"K말�5���X��m�N+zV��v-ڵj��m�2�hl�u%�9w~[n!�o�!�MY2++��A�	UŹ�~Q�������~		�EQb�i�MC�J?j�$<�J��41д�%D!��}hH4Y7�Jf��qp-���f����Hf�X.>�<}��~ V��ϼ����l=�4�\,),e(��#��L66d��#Ul~ɺ�!�<kT46c3�������\��(������_��$Y��)�^��������d� Sm�� ;Le��Wz��i(5��]�4���hD�E����x��$�˙5B�"A HH_�ܡ��I*�`��+����^���0>b4�D)��� ��c���1*����։���BH]5D���D:�fDc���ç�@�9w �6��/��l��NKw@?�x�)Ā1iH��C�s� ��\�YZ��ѐd-c�ݹ��X�m<�C�9Zk�����gF���hA�Q�B=�K5{m��ӎ�uN=��Ő��{BP���8ٙI6�M����^&��]
$��&�z��&q�9;��s��G��ޑ}Eu��n�Uq�cԮ����b)�d���o����xMjt�;����l�M�{�mSŨ����ʘ*�Jccι��Zgލm�|b{1;l�i{�:tP����6��bVΨ�29Tk�u�y�˲92�ل	�S7U�	(�o؞N	F	"i�>�D^d#����(´T�����zy�ܧ��T�R\<��
�ЈU%ǒ��	��0*�/�LR0?�nN8��o�"���#����c�M�"���R���M���-�p�	{F�����%��6*'\�Y�����r��c�C�1�D�kOV5>]���ۗ�Y[g�"�;�p�o��ݎ%ή�i�|���>�z��F��Xӄ��FО�[Gm3S�Tm���a.	�Jl�ð������SO1��ICa2Q���6��H.'��az�=�{�!{�^���#!���V,�e�Ҙ�[e�.#h�sG���zyw��j��-�g�Hn��g�`���CȰOlR?�F�T1�ni�aJiϷ�ʵQb������^�'CG����O6�ov�1	��f�ַ�sִ��T�QP��H3��GE���<��{O��4�@�:Ŷ��� ��r�ң?�������Q0J�"�I��=N3��{4�DR�Ęyf����R��!��8�Ѷk���*��2s���nl�&K
�����;��^�~"x��Qh�!⺦��dE��s�6&C$NK|�uC�TT(!sk�zT�TD��0a<1�X�x��G����*�^�t��q6U�]� E������F�	XLq$A '��Y���Y�10��
��C߰g�
��s����	��3d���MT�.��(U]#SCoy�beiT�`�h���(��A�`"!���W~����g��߇���e��#�_|��1D��Ƚڞo�(sE�����V5Bb3��Ȼ�'e��-W{����S�H�1E���X�΄�
��TnDh���PG�+L��vY�}�j,��FD(��4D��I��b��Ʉ�h@>,8{�<���Vn��z���/�Te�OW��d����;�'�QLT�u3cc6e9��M�R�m�X� A���t\��zv�,M�T���~� _iڞ_�hk0>`*O��A�I,j�bC�=&7H֖��l�C�e�:��`�������1������zwn�R]EڶM���̨ �	&���sѨԍO1QK<2�(��Q�<�;�d�Y�F�9�׊4��X�w�H E�8b{=��a���j�$� ���bӠ>U7�x��Ȳ��={���˨|ì��; �|5L;gߎ�v]�Ι�O��Uw~z'�6�U�� 7�G��%�yk�|�j�O'�����R��T�^7�Uɶo�C (��dy���4x�mm��̤j����bmj��fJ&	�o���j����Ά.^D=�(CX�{���:���-�OP%�m�}��rȊ��lpb�"̦c��3\^F�^d9+���Y�����&��H(.��e�W�GXn�T�Ȣ.e>|�����rg��"k!"�m�y��k�)�%�*z*U�(�o�94ϩ�030�qhW3Z	MK0}\������CFˋR߬eǪ����>lX�̦3�S��$b���Na��N�~+
ѳ�Y�Ѻ�6��q,ڂBO�=1ЏJO��
=g�L�쨗t�/;���u$�ź�p^�x���<��,��� �98�ƣU��@��-3��^0֠����=������ ��v��\[���Թ�n��ж',v�kqm{'�
�="�#�i�[��r~W�������G�ݮ�79v�W�6�i��m@ӥ��oHi�6Z��DU+��� x���r´�q1���A6K=��{f�)US�Y�@��Z�LM@�0��v�޴Y�pi�:ﺥR�������s�"T�3�kf��
�Yn�֢b���q]1�z�!01�Eox�x�9v�[�V%O=���"�ٌY]1�x��eL���lL�y���
���Д%ԞCa��)\R��LFa�m�j��eXB,g���KԆIV�J�b��4`��g�I���,.,�w���8c���h���7�yEl�Qg ����]v�c�ӯ�"���\�nޚM>|����,zLWRWi3s��lz����	�"4�>uQ��P	Lbd��جj��?��?{WWٳo?�++�+d�=D��	US�2�N�'T��Z���0�<�-׏Y[[#����p���op�[X����Uh]�ˊZ��|@��t:��x����.�P#FQXT�B0�ɰ6o�*�D0Q��iu���2V����C�t0�n*&iv;�8��c���:�I]�,i��f��np�ݽ;��38�%Pb�}�i�'�Nr��ͪ[��]�ֹv�ɼ�����J�
49i1��<!�[�2"�(���~l�$��]ޥE:�^��dv���������uy-篯�����/M�`�dL���Ș4�{ژ2�(h��&��5��M�,��"��[@u]�J�3�&v5���s����O�;��;�VFWS�N�`I�b��3�xk���84T��0���o��J&eEu���d�!6C�#IQ�@��cm�`��z��3�hy�ba��Y�`qy��fJm�g��]�E�ll2��b{}���p���r�U��,�=�Ұ`�X40�Ȋu�iI��E�jJVj1�Ä�T��MM3+Y荨M` ���T�.������`��_�Ư�~�So���k`��k�?��ϥ���ɼ'Ӱb�+�3W�!�Z�̈́�ѺN
A-�F����(�vlh����4YF\Zf�.N�����߻�=G�p�ד-.�-,�����<��3����g%�gSj�0�Lڌ<�<D��B�1�L��0�c�ea8di���`��pD�9V�]M`���xc�r{�l�<.�H�@�J��c_���",ˢ*��3��%Q�Fɍ%o3Hѐ��(Յ���s0������5M>���v�k�jJ5�f�z���$�TRK;��fWz�Nyz�ۙt +z�:;'!����Mԣs�W�w�rK�{GРDBv����s�U|�� )�p�s�:[��k�(��]9xg�`�k�n�q�՚c�����^"!;���]��t�#�S)=�	kS���x���,f��WH3nQ�Je!/ ��JҬ���:���`h~�D�,s�tm��<��N�ޭ��8�$�"�<��v:t.�}Hlvb��@�#�����chKꆍ�J��bs<&�a��C�:�+�lmOY[���B����^z�!fi�{Tu��os��Y�@^ψ�	=�9������ X1,�ٷw/�W\͕��2��gsc��Oq⥗9w�$g�sfs�3��|�,rF�0���l��$*
ָ�1`��PO+F�,d92��57������U�UU��s>���o_v꯲��5l�ȱ��V��W�gm���^�w�)hbׂ4lb��TU5�GO�3�lG�n�J�圬jN�j��"���v�{�m,]}���<~�'^x��|���ϱ�5fk{��t��$2U��:�*I��Y��DSZ�����@�,��6װ�F��y���e��;�b1 -����u�7S�7y�g��1#��T�l�f�B�v��e;s�$�\׬���8YF?sbɬ��Hl{��-�"�\�}Ee�s@�e?�o?�DV,��3�`�Ҍ��~�	�w�3����I���9��{v��]���'�5	���v�����}������Ϸ�,�,:E��V�����I�'���"��!�[f�T�m�'k�||�\��_��U����ܢ�B|�Yw^��NB�Y
T�1�rJ���Ν�gM����h"?�9�E�4��4M[\K=tθ�^�׎i��̈�;t�T�kQTS�E�D�L�lG�3�Fb��	[�n�2�m�T�Q�'c��	���G�p�-��.�ǜ�L��S�&�x� �������k?��Z1++Ɠ1M����E�������\QPH:�
�(\���"{��p��!�=ƕG�ྷ�Ko������<��c<��cl�K�&�8�:��7���7X�5n���
O��&[2���N+j��.��k�N���-}�_��ϢT�D�ɘlq�M�W?���I�����_�Ez�PT5�r&ú�2���տy���ps��Z���ɩ&3�"j���B?�� ���4�X��m���؆����w��;�d�0���|����#s����	����קp�tJ�S�T��
�<��Ysi�*#�������$dj�!�G��bqQ���3����=��\�����S�?q�rs�*hf�o����c�1쫄����YFY�P,JJ���X��Z��m�׹%�O���f~�c"lFe�B-�;Ωc�c\��o(���Y�b����q��E@M��T�	����$��'(�L��9��@���vb	Ӗ�Ud^�9���m�䔍5��޲�S�ZQ��m�8��"h{�B*�w�:�CZ��+i:�7���:}W�>�j�J��D�'$�B��Db�(ubN;{���W��şq��>!�w��5Dl�PUʺ�ǈ��l��v4Ѷ�o1�,sz��I"������^s9b�+�M��:�u�B]U�!2	�M�$*��L��|5c�*i�#_X�?r��1.�o�1����#C��g��%��*�Ϟck{��g��*M���uL�YBK��@��b-�&0h�K&VEQE��́�ը�>{��ppu�{n��o���W������O��7�ͅ��'�,9�-p���h��z��)�I�W%+zd�!FD���Q&�)�&ۜ�}������f�[uf�$ϒ��������7|O�,����;�	�i�<0�}|�7�%��O&c]B�����6bSUf���p@���%&.�|�p�*9t�ͼ��{Y��j.L���C?���.�?�,�	&�ٞL�{���i���4�]K�b�eES d�eJE��捀�I\ݚ��$zJ$,P8˸.�9�ha��蹰y�'Ο���/��+��cW�r��g�1�p�����7	��6�ͺf���hΐ�(�RX���^��58�ȏ��X��nI5v�C�mW�J;5 �k>�'4	
�B	V�>��P�	�=�=|ì��<�Y���xz�6�N�m潫cj1;D���l6g��n�a�3��3������V#Up�N�a�6���1�M�>�5߮�1-)PW~���{#N����ۮ�(m�׮�-1�H��N���#��O22_%�]=ni�5�SU�o^R+L��gZ@�I�y�&���b�]e}u�hw�BS�c0�Èཧ
�a}{��|�`�[6�g����f3�UV�)��Ξ���e��C��t���[M�v]Q�xU��>�9�F�l�X�`8DUϦ�*D"�٩F��xI�'�	��ل��-�|�,��a;4��:ɳ�_�?|��=\w���~�m�x�M���0����_�/|�!~p�,{9�����V����'��l���J&��t�Noefk,̖�r������bO;k)��]�K�]��w�?��_��2���Yl�[��o�>v�����'��e�C��lO&Մ�	KW���ú.*�M��k9z��8zϞ<�|��|�����G�52\Z�d
�ʒ��Mٰ���4�h�@��Ǎz�uh�1�^EU|ܑZ��>ej�2ω��J%9#%Eڪ��x$*΀3+B������H�7\⊽8���R�����ƅ�T�1�)	u�T5EP",ò1,),j�`�J�3P��������� ��;/�x��I�퍘�j��P�[�&C�S�w��ѿ��0�]Qi�/B�$�)�<5��qi�L��1[�T�|;:��Iĺ�\��_�=����e�
��Urh:b�҄��c�4���Dg"*q�t�x
��(GR�њ�D��z{>?��'����f~T����x@$&����Gs��%��x��O}�?���Z}?�D�6� ��ke�4���7�c"i�E�5�-"%������w�A�O��"#lO�l�J&)5�9#�+g�Uf%����x������ɩ�g�T5�`�p�
�zNm�qzk��	<�r Z����(�mPV))��o;a�6�����>�^GL�������O�g�$V;1������oe[��0����z�[���۹�Ʒ"���扯~���YV�!�XuaV1=�������Mr���{��M.n�SŨg���A�����s�"oƣ�����O���'��r���
gq����<���Mt��u��%�B�J4eY3���B�o�ѾػȉjʉYž���m�����y��o�-���y���H�8��+0�Q5	�F�#����},}���e��@M���&��1�	Q���4b�E5���OFa�Y�֣'�brKV��/��{9��b��K��)�,Q!+��B/p��Y?w��.�a�r��}��z�l���Ӭ�=�,&�P��3�>�cĈ�fh���:
3�J��6�횦�|�-��لo�<�B�g*�!b}`<'��k����>XYFM
yf��vNEZ�l!R��M����n墦�{	m��I{~��Fh|z��Du�FЌ��Q�t<cR��C�&$VB��90kW������E�d]�c��i�s\T�3��O��̣��#"�	��9b�ݥ��}+�y���U�v�M�ޓ��-�a*o�������u�c�ͣ�o�c`\���cg(�0��b��k��p�-�����e�/��xk�8�L�.VlWS6gS*�f�S�PǐT��	�r�a��A��Aiꆢ�c���p0��h��PM��*��MŴ,�MK�&�K�;b�:�t/K�V��ѐ���[aa踸~��|�<��Ǹ����y�=���;���w�ͳ��./��&,�,��EN�6��Nm�*�ل�~���1���GWUM��\��r�g��CQ�(�sO�gb�3����'~���b��ecF^�L��Ǟ`�~V�U?�0����e���F�0](��K�e��	q�
���x�<�4��ܗ���Oq�☦�D_�wq�1�������l2���C��#��
&[T���������Y]�,K��!�3ơ-��T0u��<	�QLa-/��yrP��Pe6�&<@]'Н*�q�2P���,b92Zb�`����E6�b]a�^����%1�X�j^���Y�6e�1bb�������;��ֹ*�(vN:�J{�HFאU���B�Đ��r�|��y��CGx��_�n{+:,h��\�D���ib��ʕ�,2�M�%iv\1ږ-S�f��L��w�k�1iuv�bZ��	@���ۆ���d��8C7f?�r7	q]�1����g�L][gCD����m��<wg��t��Mw��Wm&�~wwY��i��m$��i�QԤr{jE�s��;���~�S��\�9c�����%��eѻ�u���T[&���������,#�izՑD��x	���A�*NK�$BIs�U��7\���	:�qn<�������\����E��N����5B4�_.�f����ؤ�}QP������i�C�2�F	�RّM�B�k,EQбf.#ϲt-�=��\J&��ǔU���S՞&4�� ��r��,����d���A���e�:|��w��6r	<��/�����	�[�\��,2}�E��ֲ9�$��={��Zx�Y����\���z��M�"4�>q�*�s���^��5��zk�^��R�d!,��|<���X;5Ö&6�S�z���5�0W#./Q��ʞe���.֬�S��*���Os��y��h0��0�l2o��B,G�p��r��!�<������x���:s��,�b�c��P�&m*u]����-�e�׷��jMA\b8��ͭ	�$1�Y�p8��P��|C��d<'�&GR���򈋳���s8tp+f	��T��d�!�d�vUQ�2aC�5߰"�d�u9��F&��3��4"�:Qm{�
�!����Y�v:��^�ˉ�zj���'�?aՂ^<͉?�7�w�Xꖡ�D^R$�7O
��H�gm�1�$�s����&�"�cr��k�K����Ђѻ�sHzM�tm��Gh�Ĵg��'�<C�	���D!�-��xfhlb\kk&�����M��� �Sד����;�`Z>xLD5�x�X���K���H@���� 㪦?��X�з�zF8s�_�
����&,�������ut������&��3j���鞣^^��w����7�B���3���P�t���8 ��$ j�[���D�*yA�����)MCUd����,g6�)Mνx?������x�G|���Ő��'e�~�ٺdC�邆��g��F��d�b��ib�VI8��x�Cak���I����T�s�����c��C�Y�`�B�XL��_��5��g=rg)g%��}+�(�"p~��{��=�o���}�W����?��}�e�������������J6����8d
�o��|ع�hf�_�0���m�g�.g�����~�\@&[��,��]M5�����vCȤ؞�4�r��&5۱f߾��d��+�#����W_C3Z�;=���MN^Xcmc�Q�"�)��l��3�l�+W=�o���n���`����?��<��O��,.�V(������$'���W�{e1&E0����9�o�~�e�kb���(
�5-����ˉ�91g��uE�<'z�ͫ{�~��ƩS�x��~B�.ghU�`�}�`�GF�g��ql��P<��S���$�av���*��$ܭ��Sے����i)C�r+�w4J4���4Gm�E�8;葽�|�����@o���!m[BL��(N +-;[Ⅷ-��4_��y�u�%żZ�B&6�6��v*@S	��#��M�"1��B+s�|5Nhe���x%V�>��1Ks�F ��_�t�M��L�4>�e�yùm������MC��lWۤCB[��؀R*�������@��2{�9���\�ރ,^�`��aXֈD���tH �Ԛ�͚�kd�j�d���~+o��z� ��Ǘ3�C�r�$g����}�Q]3���L*U[�u�
u����i�fT&�e��f/�TS�tp����̹3|�/�����0"��e�F�0�2B%�f3#Zig���΁+:Z��!��:w�CR�b�O�Zu+B�gmpo[����'֚yy>��1��t������`��pi���"�7Z��
^<�2�7�x�
>�p��Gy����������ڥE�	�O?k�,�0�hɋ!��|�������L��O=�Ci2�o�������5��Ё���_��%v{�a9[����=��o)����,�����t���[���WP�{�#G\y�}��R�O����7���MVb4Z�5E�S/�`����e��N�~�mh��or��9�~�i.\��2l�RZZ�'�q3wĝ��8�;}���彂#Y�Q��|�M۲[w,�}*ωPV5��{�gyF��8c����E��9�h����{3ǕC������=~����D�)��Y��J��`9���1b5���>{�N�m+`Ρݖ��$O�4�a~�ġ����uhi���y��hE��`A2��9k8S8�k���λ9���Ɏ^����� à 6K$9! ��&�!�~��Ͱ�	J�l�C���Ӵ�9�>/�X�:Z�'�kO�8mI˻����~�a^_!a3B�Ɠ~��f'ז�ηҚ�j-OyL�pF�.�6�Ӄ�QX�K̺�.�b��w��A�@M��j������|���gY�s@aaV�j��ƌM�޽M�����-5\\=���q�-�Q9��0''�u��"��\���M�x���[?x���a�DL^w��|�\X�b#U�36��89�fS��;���w��g^~��|�W�1XY���6����H�����uS�m�>}�i]#Bq��:�M��!�$�u�'t-*�	J�	�!w�<�Ӿ@HǗ�wo��Y�f�>�8��{�P75�ɔ��Q�=���b�g�\�ַ�gu/O>�$�|��޻�����u�m3���w\|�q��
g=��'Y{��M�D��!Ő'�Ӳ��Ơ�����I��++������?�������_k��O~�,��(�3�X���n������llbs�Zl--п�j���[��,^u=��x��g�7��<�,G����Y�xVRמ͵Ν8Ũ�����]w�AS�x���x��l�S��n�^���X�Ռ �3���KD#:�FU����V%�c.�$#��>1�Dm	��b���F*�E�4~���x�4�U�hqč7^�h�@��΋�=�b��#�?�
<���ʒ0��6q�){�a�f,",F8�,�9}��E�֞<���۞���,I^ڢ�����;Z����	.s�t�B0	�o�4,��3�kְ�Ϙ./Q\{-�o��՛ߊ��
���_��g-M��'U\���$YJ�(�@,�v�������6�j<4>�w�	�n�ܡ�c��z�V��8Dӽ'D�$�W���o�����R������i�=6�Gb�uݤ�f�I�{w���e��b�F�C�kR�{>�i�����ŋ��x��K/q���ƞ=�RS1�K�MCOH�w���p�CG$��`�E\R3;W�=��_�E���Ø�o����Gcdsk�ǿ�U&/p��g/�ѧ��ǚ
�`o`ҔlMfL|d���ZC=��̅L3���ˡCGy��'y��9�_s��x���8�v�&Ϩ�ej6gS��hi)�{HR�u+���V4ۜ�s���XO�1]Ʈ-B_ ��sG���:����g-�^c��SPA�4"����>�@���Uʹ*�:�9���Z�~�}�r�-�<y����׉M�b����^u����O|���8R��N��ԣ��[c��Y��������Y��W��OfY�� w`Ͱ�o���#v��}�k�C��������%��1�!|�4�| c��$��y_���dx����}�6��︓���?����׾�s�Or˝wr��w���|��/�`��&*���>���e/Ͻ�Ͻ�gN�f�=%6����963��d_*[�q�Ͷ��36Ɛ��%�����0w֩t����꺞;t��ń�N�1v�?���ጾ�|.�_�{?�o}�[���[�{�/>�4_{�1�;t��7������R%��F#e�o*J� /0�/��;z��\��g�i�J��ٶ����?�^f�@�<d�+�����Xӫ�z,���sl�8���|���a���2���b�M7B�ȑΡB�-W��U�
�x�2�!�ʊ�C�Μx�,Éг9�uĺ�)�t��UESթ����3@��
H��<>l�a}4�x�L�d����Ф M�bMFY�̦3ʺƇ� j|�ٽ��ľ���Qi����k!;��W�+?j
$Z�<u����+ U���6�[�_>��>Bo{�bh8P���cCҷG=j"���33/A3p���sq��П�[?���_��ϱ������������7������d7=���'��J�!#L�s�i�PΘA����k������������p�;����>�v���*+<�e.�oa3�B;���������{�[Oʜ;j�v   IDAT���Akj��-I\�8�礻�#2i�~ަ�@�:���h�o�m�em �(R�.�-�>�����9~�$�Μ��-��?s߻����ͩ�'��?���}���x��������|�K��	�^s%{Ey��G8}q��͔��^FEqt{V��0�	F�3uи=��~��w�����	M�k��?�w����ЋQ�͆��n��lqo4Uɴ'L�dW��mw���>��C�����ԟ�o}������?���'���d{c������s��aV�~��N�����	XC��UM�T�"g{��d6k�R�����^*���������y���i�<�i���UU]:���+�#���fi�@_�U����@�ǟ|�������?��_���=�ˏ=I�#ý���<{�m=�84��!�G��h�,�l7��6�.S�P�DdN���W�\�:�=�S��m���]��y���mQ e�HR[�>ҏ�O�P�@SO�=�ճO��QdSky2�T5���j���o��ۛlmm���@�eq���0ڻL=/<�RW����,.�g���~6�b�[�Qpb�<���|�2�"B4�`Ӧf}{�2���Q�oq�gq!�G�ɔ�����PMcOM�����g��р�:�,g�٤�݂���x�g�@Pi	�b�x$�?Bi�o�}��X#du`�:����5�t{#��g��@4i
C��*6�a��m
zS���=��~f����3l2��=u�$g_~�Y�/S]��f�h�J���cj���MÖ3�YF4��N�cx� ����.�S���~�Qo�kn�����гϱe��*cWpq��v��%}�ƚ��T�Ǌ��Ƙ�����䈭��K����������H��$L[�`1�1�ڌ�m���iK/�R���mG#%�VF�@(����},���l^8��>�</��,����p#��u������?�3_��{7o}߇9��üt�$���V9���2��,Œk����_�~�m�Ws���l4�G��0�����?�g��	<�Ϟ��s������s,���t�0���e�7�6��;ox���a�	��>����}�D��,��=��6���}������x�F#�����׿��a��^�z�ٷ���~��?����(�dL�+--R�%[�	M�@&0�=uE/��Ś��4w
��<R�#�2�<Oz��SV%Җ�c�Xk�}�$�E�:w��.�|�$�N+<����{����+�M��x�S��h���ۿ���^��GE���׌C��gZU��J��(�g��&� >@���sh��i�씾%M�ԗ��ժ�֣�r{#bb�UyKT�ɛ�ֹt�c�<o
u�8K0f"�Z����z�M��B4���hmAwK���ǚ�9(,kՌi�ɢ��ܼ��"gu�>��		�[2+�%_�ܔdF��b�!4h�I��))} b��W6����Ra�,��j�,�AA���,a&43L
GR�MB!*$ �5i��7��9���	�6G�[@���ӕ����}1��<G��szVm����l�P�d6ipC
����O��'G��Ǐ��4��i!�߁pn��K�Q�[��wqm��+����o=A}q���A��e�e�<x+\����Jƪ�^��ڳ�>f����_������C�\�uo��G�~��έs�-��&5'��y�ɧP#��Y$s�j��d�E�k�X\�&S����~>h�%ϲ6PJm6��XJ2���W}�W�ˡ'V<�Z�_�*����+�,k�F�hP~���g	g�*��}I}Mn��#ʪb:���y�Q�_����{��>�k���>�q��}|�+_�S��2��N�����޷9�ҳ8v�c�����L�j�Ք�E︊�\�.1|5z�i��,�7�~쯕C�����c����Ç)�����m�4[�w�ęw��? �QM���)�?�\5��>z���z/�<�g?�YL���_�8��z�=���?���Ʒ���_]���ceq���kl��c��c�L�jܰ��DP�U�Zl^P6�e9u0��p��C�w��.K/˒�(�<FM�-">�2�vc�znЕ�d~��2��1���D+�'+�^��d�6��7�Y��O�+�v���{����r�ʫx���s��g���{8��Ӝ}�9�:�u\(+B�Uк�(K�b��:��䭃�*��7�:��� �:��i�V���>Si7�T�5mq�'�,�ڧT3�IekW�2��E 6X����?{���ٙ�wb�'����O刪BΡ@�f�MQ�1�"(�$Rcό�/{ֲg4�4J�%Q��83����h42P�@�N>o��	���s��<�!m�{�B�:u�����}]��^���0n�΢hpX�ʒ�C�H`��z��c&�E 7R�Rb����Y/���gf��c�
�C)~��!��`~@�B�D�I�H\,�)�XI� �EOj�I:y�3P��
���uS�`�-�������d�\'�v�v�o�>|?w�iJ~���O�X?�a��
���4T��o|�U�@���"@����.�`��-Vx�!��I�h)y��65�d�p���e�{�d����i�$	TKjc<��Xk�ZQ )�բ!����?��\�|��x�Ǟx������t��M���#�4I��9D3�v�6W��$r�Xj��qZ,QR���cvz1-0�E��=N"�4�����i���uإ�ɝ�@�!� D�ֺ}�{���i)Ňv��"��h�V�EG����T(�����`R��^�Ʒ��x�~�/���a>�������zy�I����\�4W���G�����e|c�Bo�j���y���oԊ���J�џ]�̟����RT��//������/��u����3�-L��A#��jf�����#�)s$�r��m�}�{�ٳ�ǟ~��Ǐq��W��_����ib!���s��A�8a��
���q�!�t�mͤ14ւL��'Ja�����8��<I�ɓ8<�ړ���JVUi;����v�n��|G��g�~���K٢E%*�(-ѭm�{GU�h�QyNU��ڐ�9�l�m��/��S��/�W�z����g�������^��k�@���:`'UD�ŬWI]�0���C��ꨜTu�EI��u]�q{�4NX��GEW4�1 !�� A��~GX־��;�;#�69KȰ��'4>�z�RU����z:"�N�p������t�5�EHŲ�l���Txb~Z�exh��A9��-2�ȉ����v7�~NJ�@X�wES�T^��x9.�$O2�������(��2��=�S�=�y*_ǂLš�߮@v����G��������|�����v^���M��1.��"��w��v���R9&Wg����y�;S�`F#��~�h�<����8��d�^�@{j3��$É�n<)Y-**��,+��>��?����y�����A������ܜ��nz�9^|�Mֶ�(�2??��+�7�0ń\�� !R:�ɴ�I������.��»�>jm�ܷ�v�ڊ�RA|��zp������ +ex>���N>����J�O��y�[�V�[�b��{�N���EXG,�x̷��*E��_�a�8q�����(6VYN8��'�m���ٳ������ߤj&�Q�����ʛo9�|�F6*K��_����?������G��3S�����4BJ�NN��	)������ԏ�^��>{A�
�
F���`��ǉ�8Jџ!�_��W�v�<�qN�wY�p��3��_��~����d�޽diƍ7)�	����� a�T�.`%��$�gh�5gƵ�+R�d�󬪊8�w;m��n�����j}�xWU���᭵��`�����?��UE;ﰵ���Y������)Bh�ń�[�8�M�\Xd�S~�_�*�R�����?t�O��_�;���LWV8���\�S��=K4;�hk��(�y�D����5��$b��>�|(�η�mh�b�QQpqs�A�3H���A^;��#۱�oR��phǿ+ڽ�E@��D��ݥ�M �x('ClS��1�z3�����o^��
-"
��1�n<Ff9�w���V���T�����"@Y�r*���$Jb��S���;Lm1�!�$�S�8��˱.�'IDUMY68'0�`RtbH�4�i�������~l_���]���>X��9��r���n�/ي� Hp(񟿳�j�N��CD�U�]]%ۻHt`�-Qb$ܺx��������1������ΰ��Q��T�o`q��fU�nU��Z�Tq��O>����r��-�=���W^$;��/���B��W���[7I��N���&�h�)'��"�3�wj���uUQW�n7��)G��q*	EV����t����8�.�"����M˺�Y�������vRbm�h:��D*�1QgmX�(B��F�*�YFYVHono��g��x�͏�؏s�S�q�]4�Aξu��Wnp�'>�ŷ_�օ�8~�({K����[�&^�Օ���q�M��Y����n�3SлY�Ԓt�'N�ě����#?e����|U�K�5e7a8���������3{���e.]����Nr߃��}��g���ϸ|�"���N0�es����m��"�>e:�=��1��㰍A�!%��;B����>;� �63�> ��:e�5�γP�)^���x:�����;�� �0M�a�[
�l�I<��ᝧ���h,�s�t�9����˰���o�/��Or��w���;���S5��
c��1�A*��"�1.�?��[���[숮ڐ���+!$�~��FDE�(
�ip���L�0
V����C_�S��yjN8-�ƅXai���m��$�:Vl`i�0����Bc�%MU���')*M)VW�LC�D�FM�U��a]�[	e�V�mgw�~A7 E �i�Qq����p%<�[Ĥ�Z
G�%���N�T9Q�VUQ�T�DY:Q��{�t�J��q�K�~%�Ο9�rX��;7��⇣{�}X���g@(�)5�	�d���?s��5��gX�L7��Ӛko��^`���|����˜�����׾�\S�8���n�03������o�ɻW.���C�)�]�½��4�y���e~�7�#�/]a��EI�ꍋ���JG�$�ZyO,�sg�n<�l��;�m܎��sh��0�\+F<��Xk|܎�[a�N����;�cvĤ���Uĳ�c�� �1A����"���44��4ex�����2&u��ؤr�{����o��/���!Ds���x�׸�����������Ǒ���M�\y�]��;�%����>������������'������]&
�?�k?���4�����~I(��dv�����rx����b�����?���Pf��%n^�Ĺ�'?�y���Q������W��/��{bs��L�N��d<%��ᩚ���T
jƅ�Y��Þ�}�ɐn�mo�m*��d�l�������ʶ�3m�1u]�'���_;���X>�ew���9���L)gƠ�#Ѫ�Ǵi0MÁcG����|�?�S?���={�a���\z�4O|�3|���`{4$��b<a�:Y´�l�*�l�D�ڡ��Z)d(<�n�ቓ�=��DZ#��x��aT�r��?�(m;EQ��Љ�6�E�b<�}���PD�>�])	2B(�B	�1��>��Ѵ�Wlom2���v{�*�u� ���Z�RX��h)P>`YC�h3�[��� �����m����EJ{�zH`JcA�Y7"&BKx��⼧��t{��P��!���̈́X��2����i�#�}�������������p��|��F낝{�8^��������w�O�qA���<s���}���=ž�GY��I�8���fHþA���=n�Y6�{�}^P%EU��r��H�f�����,��t����Enmnp��'�̏�0kkk���x�՗9�����������D���[b��ց� ���Xe�2�����,����[A����3f��i�B�\fi'u]��X��,�5��ڦ}��V�(v�x<d�	��8�j-���H��J��E)A��a�e8-��ys�_�������_�������7^�+�#���g�%.�a����K����<�wq���o�n�	r�����o�S���NQ�3Q�;i�����<yډ���hn��nU�>�ZS�S�l����d�(g��n��p�%⾇�%�T��ܕ�����Μ?G��+�qr�����j*SSC�-��8���xM!��y���?܃*
����<��t:t�]���i�]�z�$t�]���w��Y���������x��}���,�i���m�jk�����6 �s���[ ZG(vv���M�9D4���_���?�c?A7�Y>r�b{T���#lm�cF��d8�2�eHQ��#Q�L*/Q-Qn���o��B���9�wغ���j����:�[!�Nǡ];��KҊ�`�p��Cz�[�,+Fh����ExRơ�t�n���]��@I�F���#�|�&R��#��'9�y&֣��)�Er�AЎm1G�H��DP��t�&������n��d4%��y��aR��1M]�㈬����:Mg:��uh<�
kɄD*��,��&V
d�*����ֱ[��� v��l?���o����;F�*�=�$�}{�
"��U�Dm�]ƅ�َ�l�xn}�Y�g9��O���'��C�@Z�rl]��;��8���5�5u]P
��YJ!�ğ�N�����_�����q��)~�i��u'�������3s�n��⽡��8�uYc�8AiI�Gy�֊(
�RJ!d�����h�N�,Q����EPm����;������M�U|��!�Q��U�fXc��]�]q�sAD�e�а���"$�9���E�h_uS�W$�&5�b��x�U�N����?ͱwR��#'��ʙ3lON>�1�ǎɵ���N\i���j�9�|�;����T5�!"��ss��������W��/$�?p��(�R)�n�n�/�Ts�ԟ��,ܱ����<s�C�f����y3�<��Y@�3T"bl���Gԉ�ұ��ų_����FHBjQ�$XT�J�0�m�pŴ�]��y���H�QTP��S���ݏI)���4M��-�6!�6���jت���$I��|w���Z�֡��2���-uζ�T>�5�RX��GGq�w����	�6x��*nO��<M��Q[�h,Ѵ�'�Y@׆o�ޗX�g���q���w����6���~�i�~�J	��ත�I�aG�t�.��8q�Qi�vm�.+*r����1�H�H�7Ex��S�Sx�0�)7�,�4_����ol����T��`��%U1U5Y��x2�Ơ��FkV&�v�qBm2)�a
�fR���{
�8K�U��0�CV��8�*�c=�jX�*�	�7$y��N�k�l�"��RXoQ�bn����1p��y�.
�����8�J�y�hf���6��U����kj�������k�}��Ϩ��mm�ԙAF	M3<{%Ѡ;1�VAO&x�(�gG�<{�.�i�/!�L]��;T�)R�~g�
��3j
�&BV#-2����xO����d|UKf�UȨk�BDljɸ�ti[�#�W�E�
,�u�6�}��wޥ�#a���b}���C�	���\s��psTp�O3{�)����rϣ�2�wNG����,8�W�������_dfУ�
�67��
c��HWA�n���Z�u�>,�Y�*F�1���6��ZK�i���	 B`�5�"DBGZP���T`e��Ԋ4͐���%R�:�i�R��Y��M��焷��,�TX�>Bi��J8��(m-�m޺u)�Rc�EO���^�RӺaR5���i:��Gs���#ͻ:q�[�/�K��z蓜���E��q�M��{�B�\�I/UμД�q[[�C/��T�Ο���/�����T���͒���>�-����K���:}�1ň����>�<zѝ�������;3�*�x4�w~�?��g���zR�I]c_ckD�z9�#�"��5 t`s��"�D :(%��zk��1��Ӱ���p�,��ӌ�0�e�qL���u���XKp��X�5X[�l�pcl���h%H���$M����pBP5'$Y��a��5c\;���	�m0h�H�m-UQTtzpriWo\��~�7ٷ���{��8������(g9p�8׬�y�hkdaj�%Rt� (���J�ހΩ����,&�0�x�[7�����LE�5B� JQS�9��� ��vH|��o|���[��,C=�̺����D�5֮��g*b7�")X�$�G&�5��r�sK�X�v��4�Ǜ��✩�h�Y��N�.3�r��{X�Lx套����V���CQ�\)�Vh�)M� *����D.�l��k�1Kҡ|8�T�)�a����8�©YF׮re�
*�ȼcfy/q9b�ڠ�DU�D��İq�2i)P�"�q�P��8I�(
+����<��;�o�KRT�i�@�8��\�Ҩ*̆\1�۽.��C��3�Նҗ4B�TFDN�6���:�RѭjzJ��(	�"qNRuz�w� ���`I�!�#���N�nl�K�2f�*��U�)�Ք,�IbMO
��)���Xu�e���������F6;`�w�|0�w�Mw0@D1_��Wx�;��YGQ�LF#��)��� ��Y�*F)G'N���x�������iQ d���MEEdi���Aɘ$���#�C+I��XS!�xBdLS�<�&���]����U�Ƚ=�{�Q���a��А&)I�n�9��q�i9��5���j�c^���%Y;��DB3�:hQ�DM�ux�͏���қ��;�s��In�;Ϟ�9��g_��!���
��t��X�����Vc�y[���DY¯�7������?�2�'v}��?���CkM��ӝ���SR��م�c�_z]\��}�TY��G%��~��^|����F��=i����[|홯�v�6y���3C���µ�m��XG��}������Z��6�H�V��p��Z���XEA}m�� �Ly���:�����0�9��$@b�n��IM%���i�!U@�fyN���8�t:�,K�Э�Z�$�9.Z�T����4R�0zkF�juJ����tB�ץ��������I�{y�~��#{����L[&�.W�S��F"Æi�0�{4�ce�&�ޡ�����D������=˛��T��yQU�2��i��F�����C$2	QE��p�{�&��R���˿�3ȣǠ�B�]�����W�8{����s3Q���?�S�C'!N��"�ϰ}���,l8���!_�Z�`���~��G�����>���4�?��xo��l��7�}���x��V�/�P��T���hL''�§��s3���_�MJ�`;J"����Q�����4ّ����y�_�S�ḇ���!�L�����:��1���~賬}p����,�	��DMIJ� %b���|�t>�4NJn���sc�N�FW\�r-"��"���0��=��D����j�Y�S����Xy����+誠k-V�o�I��El�,���/0���ƀ�rf�&���B1�H/��[k���w����b1�Bk��pc:溙�:�ZP˔���-� 9z�N��8y���{^|�E��~����uTEȦY��Y��oO'�MM�ۥҚ8MI����n�dY�)!���-�Q+E�5UY�45D�Pk�(�wZk�$���tL�e(�GA�+�
��NG
�4t'�Б���02ߡ�y�1�B'D-�	Z;]���;H!���uL�gX��a����y���Ӕ��ٿB�et���p�9xh/s��1�q��w�ĭ^���\���ٽ�o�/���S�x����_�~���F)��>�=ݘ��<i�)e����O��0�����#�,�y'ݻ�=�an���"JYܳ���捛��o��[[t�[7���]�G��
����A�Б"��4�D�&�4Q���HK�V�G�@��[��ئ���F��	Q3?Ȉ� h �'���v�Xk�F4U��`���)�����M�
i<�5u��R"DI��A�4��O]�v���B��C�xo)�*䍋@-kLMUt:s3�N��o��������@.�ac�Bq��=�������
����֌�a�,�c�e��
y� ff�$�X�}���]��7�A�H)�Y
!��$ɑ#t~��0����K�tLz�gVx�H�Ծam�&K�?�5�v�s3,�u���k̸�
Vf#�}��<@��0-I���K�8�Զ��Ō����u�'~����q�����H�v�cQ�I����}fￋ����<�y�)A;��R�1��&ǐ8@��Ә��d��P	^5h-ip�R1s�靧P3�>N��g�<�
�U�6�����"�3lY�⁃����~�ynlY�#t�<C;��R��b�f�G��)��Hg�}�)����r�a,i��q�"��,j�O�6��0l�Ozσ�{�����DM��cL�1^����/0���p������>��M�<�k����JF2af~r���*�D�+Pq< ����m�P��QL&��C'LL�Sq� �*jᢄ�b������g��]�=A��q��1K��=�n����\�|/=I���m��w�smZӄ�׵��R��2�����uwA/�N����&[����#���uHQK�]�l�A��]1��49m0�Rt;��ՀL�`��ʢh�qKӺi�R�=!�ET+����v�GF���ӄ� �t��X]'��(�c����p��>����'J"���֭[y�njG�X���`xc�Y*&�_���W���Q��nn��?��lA����QJ�utz�3Q�������7��U�lܢGD�>�<�@�iQ3,k�D�������oq��9�8��N�E�l��8N�֢DZE��*��5Lw2L����FZ)�3��AE.\�G�ID���wr:Y�R�A���V�Z�%uS��d$!E�C1)�tFE����`<�2�L�ޑ�1Ӫ����]+"�� �3H�JQ����u�Ó�)�>�!9oiLEYlnmП�a��y�޻9��<��O�տJ��'�_�����wr���w������X���i�*&�
�b���(�T:�D���q��ϰq�7/\b>���5۶��]������I*)��!jM�����-��UÅg_a����1�N��'�b���}�2u���}��w�tFSx�;�p��W)ooqbv/��&M��'l����O�({>�$,v�f�H���Ô��4�`���Z�Y��z�������l���l���}�	���qJ�&�#AV���?�znk�c�Hﻛ�o���{R뙌��J3��w�{���E���Kh4���"��/=8IƊ��� &ʉM��l|�kd�%��t��;�^��I�nl�"�N;�K�I����q��/�|�{,�	E��01lg������<|{~��l\?�捛�HO+Rb\e�^!}��lNy���&y�mM��b�F+��*խ�tdӂ.1�uT�P*�Ղ��1S�I:}�m�?r�'���<���:q'��e~�A���C�p<�[_��ϟo}�,˨�:d��6��JQx��Z���H���n�����$:F*Ȓ�H)ʢh�i��=H�f H��ij��4Α��Zjk�U����-�'"(�	��8�QR1)'S��%U���[�� �m�ӽ�A�ۮ}v,�IaLMGzA�k��i�tr�M�3�Y~���g�:���h�c��>�f��xʞ��eu<E�J��b��MUy�pf��:��L}MV���6jn�O���_ق��R�(e0�D�dJ�����O�z�^��fJMľ���<	�x[�t��i��a���o��w��S8�"��r�$j}������{L��\�_E;^`���gޘ��lj��ȓ���>�J0;7C��(�rMݠ���1ت
�{� ��;���FHP�J+S�pt;]:���a4�PV%E]�7)u]S������+Q�A�q�I�<�u�Vb�N�&'�i�B�ESQV�(�lm�1'�Y�t����'��w=�(*ΘY�CS6��^^]_'�[dXV�1��L�e�!C*4�i�Ct�O��M���8��.\�5���n`;J�}�1�$����p��8&R9�L�\Ed����!{�&��ߥ�ß�4� 9u��'���4���ǟDv��� w�(�~�u�7ϰ��9��'�±6�偿�c���'({)J8�N�ǔ�n�z�
^E��>��,>�dI���f�X�̧�����ޣi��a��-��o�sL��=J�9�F@m��R(�X�E:H�6��ٷ�G/,�.%[�|���ruX0������~��W��0����c#ZQ:��r���w�3�%���f�O�`����+��=sy�I9et��Y��3��$G��C7����\;O*�l�S��$��&��8"������{�n��v��+Wٛjb�� ���Ty�n�G��<ѐ&��1X'�A���H�ƺ�fZ���l����`⡮�B����J�Y<x�da��C�H���~��>�,�Ʉ��c�a}u�|G�g�=��/�%�i��:�}�8	��B����"���4I����U�#B2b�Xʢ��K�8�zGQ��Nw��;��Hkz�.J��� ��(��u�DRS��l]�_����[���;���� g�����,K�pG=����;)�Rc�`�����o�s��]\�{�|���D�0ǝ�\���=����Idl>��������k�-���loCo����"?��G��ן?��#[�E�I����Q��:s�'�}���t�:sB0�w?s��M�w��㪡3�D��$�X._�����ﱹ��h{Ӣ�u �Y�RmJ�c�$�A�<�� ��˶��"�H��N'C�����<K�Ә$�P-"�8��֐�xL��()��lmo�cvn%�!� !�!�pS[��>A����M�И����N�U�ԁ��(ˊXh�<�*
����7at��(4�>$�����FR55��t�]ʢ �2N9��7N�;���9t�N���s,8�p{��Ǯs��9�xL1-�	�2��(!Ȣ��1`<�Ji��Z�e�f�Ï3|�m��{�<�i��ȣ��~U�\h�UJ�2bR�fJ֔�kJn<�,���x��V�<� ���1��ߏ��b�z��k\��ߧ}��.�,�.�s����9���2�Ce�P�mp����7����^CF1w������O}x����/I��gϧ>ɕ7�Z�`�6�D� �'L���z���W0UI�c��ԱA/�"�=�7F���|���{�����y�m���X6ꊺ? :z:]�� /�b��,�l���h��cƣ�:�,?��0�8��s�q�0���g>��s70�3�fav��l�L���j<�����@ji�mD�E"<���I	Ыׯ]�̗�D�w��S�)�d������+�DY�]�&���f�/�(����\J6;�+D]!5�(��k<��C|�b�bu\rꩧ9�У|핗y��O1�w�=�h��ܸt�g��e�]���0��҈�dB'�~�Ԫ΅��AI���v;o��uC$4�4m㑠�*�m�v�(������hL���b���1��(��!�.;D�F:�#�L�dY�s%Ŵ���P%>���]�,T�" �����.w��;�k�j-�/���	�N�kU��-Y���&�4�6$J�#MQ\<�o�����/�@&)��2.f�"�s��<ɕ������?i��Eg�UWU4�zn��K������]�G����/�MD�'��H�����G>㶷����(�t�	���`�Zi���������Os��)&�]���(Nv�S��]z|��Zb��4�Z��	�T�cM��DZ��:���>�h꒢(��c���ۛ[TU�h�q;xW����*Y��f)uUs{k�s�4KI�����C�3�>MӐG	��Ia���5�bL7�ج+��[��"��4�5�h%h*��y&(Ϥ48K{X舘Ck�x2!�#Fۛ�q̝Ǐ������W��_�/~
���2��uN���4��)�d��j��	؂�f�]Ɠ)�)��ۨ%C&%^|Ӏ�0�]����+���,<�^+���'C����N������2�H�Ʌa��n��,�ď`	MՐ�]��g�&;�D����i�([cV^���7�Kۛ�8Ƨ������wC Hd%�|����1~�y+ϩ��L�e��in��>՛��������@��}�Qn��&�W^�[O�J�U��V�?w��)8��V'"��␋�5�<�(zq�l�az�=x�GOp�ӟ�/��)�kC4���g�)��*�UB�4���U��زD��u���<���\�A��i.��.3w�������2�	3^MK-1��d]�If����P�*�n�Oj��w�^�8�眽9����?x�m�R�B޺P���S(F����Z5�zBka�&#dqim\��UL�=�f:�e�v���p�������Cw{��H����+K���op��y�4�9CQ���T�{DcUU�r)��6�8�y��%�6���X���t��c��u�-
���XKcB��iF�����dLQU�6�#�E�&4ƈ���ɩ�cΞ?G��t��hHEeIc�!"nuS3-���k�wHu2�b�x�؁�Z��xL��Vxlq�6Nk��)�NG�m�"M�5���7Yܿ�Sޏ���e6Wn3���;����6����z�<�Ī��ͧ���ι�pƚf<!��f�tI��>�=��Y'A:�O��?��}��%)�c���?~���#��{ai���d݌��(�Ϟ���{�j2�T5uQ���mX���Q�Q�ҊF�$j��*���C(�5()��07;��"�׊)�tB]��E�h<b\
�ex�i��"�v�� �I��4�n��`����h�A��4��U�iNԏ)ʒXE��w�^�a4��21n2mY��k8���i�mʗkcq-$�/����"�#��f��277����������������cm����t2�5%��-�b��UM�Z�HKm�$�
#�Z��\�@�<J��4�,=�8v�K=A6�1�B#MJ"Z(L-%���������7^���	:��i�^��O?����Ր������~�x�PD��q5㪡?�(��ыb������
��8��pp&�W�\c)�R8ǭ��bm�>��<N��S���e?�	ο�ecIjˬ�1[%kϽD����,��,�__E���Ռe���Hť�~��l��K{�&̡�i֦�BRH�9D:;����}�y�M3]��l!������al��"{�&cn�~y�B���t��c�C�~�6�6��$ɐ�����n���:B��� �(�rDBC��Z�t���=��	U�x�/�Vx�1J��Q��8�3��rj�Hh�"��4���&��3l�>�9��r�~�)��Y�/]��=���Β����m�|�"/����6>��ށ���4�A�Qh
���E�-	2��g~'�.��Ra��,^�4�7�P��A��ѐ��QZS6a/.<'cdU P����;�����M��Npƒ�i�Y8�d2�ZGG0	�V��{�yN�gP����P�]1��@���?'뇰�@v$��!�)��bM7�)�����uM1�D	�q�=G�������4�	�����4{N�d���h!�ǵ�Y��-<7D�x_�^���~��������?�]HA�II�H
[���N�y+���kč%����$��AXZ�D1��DI��,4����W_fkc�~���uݞ8?FH�kK���;��n%%���qD���56�Z�#KS��y�>�~c���e��pHQ8gh���tJi=^�x�&�y�
�5y�2�&��8)�77���iBSU�1^]GZ�u�=�#��(�^����ü�����y��BE]W$I 7MC �8Z��nh��]؎q���H<eU�]�����x�;��g~�g���H�t�0[��;z���:��bˆ��D޳��D�"O�*b_c��Z����J�R�����
�����#G�l��k��$"�T����A����ƒ�cz^3�t�⭷��q��7^"g��P�%�5de��W^b��%�ǁ�筠i^h�8��Dia2�<���pO�gƃ3[d�ĕ�q�4��/|��c�����J��ȗ�R��Zz2��4��6l�X�bJo�K��8w�j��=���#0�r㥗Ho\c��i�>� �s�{q/���"����Ȗ��.� +
:��q^y"�4D.�˄�����KT[C�|��-�m��o2�o�d�&i�$�H����� ᑭ��y0b�F�S�����c�d-ɹ��s侇H�����xrT�ܛXRhIGh��0�+z@��NB,c�ڠDM&,�;r<I�0^35㦡�#J)������|�w�]`v�^zss,�ۋ�S�e�׾�Un������?�ST�)�o>T�C´�)JJt��eصc��C+��4IEY2��8[����""���d�����s�\Ԃ��݄F�5i�`���X�"��q&E��A��5Z
"����N�s��-��Ÿ�_w����90Ƣ��V��%	�s�,4�n��y�]���#�w�B�����j��CL6V�;~���g���+����Ź�翤���h��S:�G�K������VH�w��t�]� �k��7b��NWD��;D��n~1�SU���'`LMcx�Ww��4���)��:�έ8ɦ,���0.�Z���(�h�y�$ \����:�ш��5��;>�L'�ik+$����=�(B�4K��g�.Qn'�\ :��]N�4�f�$MQ2��O�^b���*����M W%�^�!�4��C666��%Mݠ� �2��Li'1��[��	A��1dI�WdQD�4L�3�ؿ�K�q��U��;�hsKK��8z�4�m��!ڥ���TxBMJk�xC�AJMc���;)��,b6K�8G]��>W/��Q�c�#0(��jF�U��Ԭ��WvR������E�ؓ�\�b�CU�D�g�1�ޫ,Ԗ�<CO
�#2I�9��1��.��	b8fV+�v�K<�2 
��1�RDՔ��|cC~{C�*�3(�0P	u]���9��=ʕo��L&l{�쑣DsKp��� ��x���mG��λ�|��$Gwsf�A�5�gؓ$Į��ph�y����)f0���"�f��-�Y0���8�:�O?A��A��;I��;�b��*D$���ת�$��k��x�Y�h�d3K����?�������^�9s�;T��� ��V�BI&�3�$���O��#$M��L.K�:5l�d�W�}�R�ʈj\�H1�k��q��)�஻�dϡ#D��{Ck^z�4�?��6H%0uM�!n�	E�;� U@���AXk�����a
�$I��d�i"�H��$IJѴcu'<�;�4CD�����%=uS�ؠ��J��"Q����?�f�U��V�=���hiɕӲ$It���H!�!RC��ǟϻ�O·P")w;y�	H�8&K��(L�qPKOQ�����ǡcG�#�����}�6�$�`�1K'����gD�]쵍��V�ec���S�n����|}�
�V��%3���*������L�4�0�� Uw��!uD=����8o�M�pk���]��Wq�P
����s�"<+Z	��e��H�R��.�Ii���dhG����n\gum-��☢�)j����	�JIM��anv6���ξ�CqK�4h%��,� �D�)�ф~��Y���E��6ٜ�dYF�f�(f�9\U�XO"�NN́�X@q���$�����6�Z�bk���ts���}�Xoq�rh�^�6�x�g��?��H�.����1�38~��[��gf(ʊ�	"�q&L ��[���7N���C��{}dm�*Ô�X�V���׿���c�8�\�w�{���4m��D�!�A������{���_g��C0�	jd4Z%���Y�ҷȮ�0g%}g�T��!pJ������6��-Ɠ���)�	Bi��XS���7e�jC�$1D:p��ئ�G�q0�u��8z�2�\�v��4��%�>q��7�@o�&m����Y}�M��,���qF5tffX<r�N�ao�s�W���@E1�.�% s���9���ч���[t��nl�Z0]_ǭ��{���'���̡�	
jOx�X�0ހw�N�{>�9��D�o�o�fTN�=?����(���G����m�D�1:��ji���� b;����4E��,��6q7;/]a��Mj��a�.�h��(�cO=��������O�ɑ�������~�Օ����	��C�U��4JPR��rj-w��)��"˲��2H��tr"��Z�j]��i''JR�EIij��q1Ź[W!O=���8����괳&L��b�%�4��H�e�Q���u&a:ҸJP�5�~7���&�(
�i���}�;�x�u46�j���#��XO�F�a�4��4�ɔ����ǟz�{Nއt�X1t���l����{X�p�ق|�=z�7?���f��n�N�yί��_����-��G���BS^b�}���.w�7��������s��73s�"�D�m�{�y�M>x�=b-�V��6Rk��S�M%eY��o�vr�5YEaU�S�5t҄���ͻ��aRLhЉʪ�5��Qؗ�]�8BJ�R���$�(:�I󔝐�(���%��ԍ��\o����F��g,���h<b4�d)��A�.�-�r�?�37?�s���-�ԤY�x4��,c2��R��d���3�SG��(D�N��d�f��^{�%�����'���0��{�����Romu���
W	l�x�qu�ßy�M���`��(��lB�b������z�z ����0��+�Aր�2k
30��w�1s�<��O�����p������I��.+��%�Y
�pe	*l�Q
��M����Ǩ�&J$Vx��h��Q/G9�L#(�+�l�����m�v7�z���ϒ,�=y���o���qw݅/V/�G�6I�e8�y�*KÚ;Oq��Anom������/bV6�h�p�CF�D�i�?q�g�͕ۼ��g98�2�c��Øs/<��#������n��1P��u��Ģr��u���rH��03����:��WO������`�"�LT䉍�+-yQ�p̕o����&z:$5�4$x�t�eI��n*&J�%צc�=�8����W8v�$�$GH�u����k�r���H��$N 
"ٲ*�"X��<ψcMQLC�Ob�(
όv���)�n�U�B)�AG	2�0MC�<�"�S�wL'Sb-IM�gH)ڮ<j�kMHđ!�-_�'�+��4&�R�`l���-,��9eQ��r������Y�Z�<'��س�J��1)��3y��&%�{�e���"|�J�d�n�"h|�I)i������?�}��9H7_�;�`v����`@������ ������C��sJ�7��7DU!�E��������W��V���gz[g�˸2(�?r�g?ji/qw%c"�����.y�7�����eE]U���hi�$���1�b�R�$�đ"�aG.}��I���t�qq��l��TU�S��ߧn�`�J"�8�u�E�<���=yY�����X�u,�/��#�pש�p�2�N��s���\�A����e	Jk�eA��E����e���<U]���t�h&#�77Q͠�ev.�P�b��c�kH��&���c�x&h%�����
��f=�mO&t{]泈c{�l�Y�����):��3��Ո��{Մ+�k��r� ���q�pF"�&rp�*���W���a��{/�.��`+�����M�z���CPj�1DbO�kb_�(1��`I�m{e��KWYy�5=� ��CH��gΠ6WɵF7�kж!)�t�������Op�;�FN*�ȽC�N	�Xs�V��}�������w �d����hd��X��'l4~� ;tǟ��{���EĠ���sl\��ReI�������9����~���n��sߣ;2��k\]ӑRg�2��_`��{P&��0I"���L��*�46�t$,�<�����딓	�(��>�༰xgZ�q���N���{�Gz�����-��G_����]\���0ɐaeQF�K`ʍ��1|���
5�U	��(� �,B�1[u�jY�![H�X��cO���y��Z^F�$����T����\�|���B���E�s�����M���$Z�&JI���,K�(����Z�¸�!���4��n�b�]���.��"O2:yp�H)[l��6 m���()�)uQ����둤)RF$:"MR�14���)Rjffg��L�c��`��M�i������=����Ύ@N*!����1� sE$e $ZC)���H���i-Jjf�9FN�t��y�O|��C'O���,�a��mf�<��s�[�3U�t�'_�l�BcUVW��W�E+̪k�dl�7o�ӫ+^��d��?3����&�M�j�Tξ�7�_'�2�ׂ�;βݱ��#1W�D�խL��V)v�R)�:=��~H[�=������t:	�
Q���qQ`�evn@��B�x��#�"&�1eQ2�(ʠvW*$�]�|��h��Xgqi	%�Ξ%Or�f���1)Jnݾ���L�cb��������L,�a0�����(g}8�6��^���y���	D#p8�<��u�'duk�I��$M(��6d����K"�3�;����7.��s�p�}g&��)�M�<�d}���<����j*捥�6��#b�M�]�d��M�~����#;z�S�q��o�\��>�rp��xS�#O�'h7��
�m�D��\F��0#���k����%�Zf�4ʐ�
� �����0|��O����#�Ơ�9��~�����U
Ӱ�v�dL!-�"�͙'{���~�<�N+b�p���!�7>�	���%=�Vl�����G���9��C@"���\~�}��a�v$���[�]����}��O`�]�������w�n";�F��J#4�`+����?��%,�q�/���"��Z�L�nf@�4KCL��	�d	3dR"�#2�lV�����9�[�Ý�e���#���;����<��ӌn=�/�Ω�&I*�VCQ��d� zՉtzv=B�A�Q�����`"a�,E�RIɨ�8~��,�;«��O<��4�A����Ϟ��oaC]�!hl&>iDO�Te�n�iB@S�H�I�& �R�9	ޙ0~O"T1m�E��p�<�Ҕ��aU+�k('%�,��QxVd9*�PJv�3k��1m'k;\o�)l]����v{8'�N&xR��L'q���~�t~;���t�N�L�%ݼK��G;SU%��B��8B��X����.*�1Mô�PiD�I���I��h�֒�.׆c^��{�ct{�(˽��U⬋�[�ٻ�ޛQN֕��1!��¹\�SV����������?�S+W���>zPܸ�n8�tN�����D�Y�-�C�	�F���`2��k�����h8j}�Q�9KQL�kP�k%J"��-H�\��Cy�u{t�}��`�g{{��h��RQ��Ɉ��-BG���{��h���v�0�Y���9y�G�z��i�������c�,,���^���>��[�����t2���qBof@S_�����#�pi�2k+�9�}��aRLI����%VWW�SC����Tj�Ry���9�樃�N��~�.F'Q`��������0�vy��i{�=�3��Л��*�\�������ٛ��$�[��iS�'$L	c��1{�ƛ�9��2��g�҈��^`�W��53"F���ۘ�Ӷ�x��'�@I,��D�a�<Ud@Y�p�@z���Z�Q�@:ւ��RӰu�6��M����#����_�8�V�x�jm����Y�:y�SO}�����	�v{�*���,{E�(�wx%@B��q�	W^}�ه?��z,?z{����-n��n:
����*j.��bvk�����:�����.��Ѵ���HS��G{���6��=�E�����"������#Y��2��e�~�^���[�5��k�SA��剦D��Z1[4�IE�ܼr���z��?�E�=x/��k7n�מT)����,�� ���$*2�JH,$�0VA�J�N4�N�5��4R���S{�mgH�ڏ�tP���X�m8{��n�B���j�֠��/�JR��q�DƵ�)�'�CSQ7�����H�c-E]��s����07C�elnnP�5J
fz�.y7'N2j���!٭i�9���H�dwޘ�������r�R�n�4M��0�JM���%}N�u'í-�R����$y�c-��%�FC����m�Au/	�����S�(�z�mw�q!�gG`�`y�]Ј�Ao��s�9�<�H��$*�����f�:��y���ijӋ-w��Zc'��Q.�J���dA���o������}r\�4��?�X�E�������C�����9{�uU!Ň���8k�2D��0�u� b��ZJ\SaC�5�N��n�L�c��!Zk�X__G+�������yF��ٍQv��A��Y�������
�ш�8���׾J����5i����r��^?}!�9��>[�C��!�`��~F�1W�]���D���z�MU�ʘ$���z!��:�h�5�8M�6j}�v7ѩ1A���4MF:

a�N�Ŕ��.���7_�O>�R
�`vn�f�����3W��#��d�Y�<�T%Y��7�ؾu���$^r��ϰ����K�~�Kpm�E�De>O2V��x/�tB�#�	�K�$ʃ�*lǂ&vxe��!|k�*��H�#
�m�Dt�G�mq�[/p����%(����89P>���:��b�O���ħN �>�xJ�ƈ�+\��WQ+k�+OV��%USBS��1�V��#�N|�~T.���{����X��YM�lM&4FP�JD6���]�Q䳳�~���׉�]T1A���T*�v?���w� �����M־�2s�E:�X��.γ`{���ɑ�,�I���9�ɧx�����A��X��;�^UE3���ppt"&�)��}w��у�����g9%#�R�Cx�kB����x*�ФY��8���@DBǔ���²|� O�K��wם4����<��a<~��i�bJ���8P��ζ��c��dB���ć�NdFʰ7�*d4x�L��$��
(�<G�K�.amp��}�<'I� uA�R�v�xR�µ��;�h;W��H��CY��	k5���G*�e���4��Xjݙ>���e2�R���=�$�R<�r:���34�txv����w�v���:��"���8@k,Ji"��C�wnlr��y��^�8��,�֖Π�8��s�[\f�v�T�{8J�~gݪ�����[>R���_��8�x�G��kkumnvd���D�K�<��-�U7�e4�����իTe�R� x�u]�g)��X���!��B5��!�BD�8�QZQ�k�8!S:�>BK�/\�Y������h��뒵�5��)I��0?O���ID�h4
���}XkY__�'���~�����>����ko������"i'����7��g>�g?�y.^�µ7�R��������
�O~�iN��2��-._<���,cf0�h8D	��ķ7g��	<��Z���܇4=)U����ǎfu��dB/�S��bd�1����.9p�(�����=�~���y�Dq�:��
Y1��3�Ҭ����s]fW6�F�B �Eh�wN�t76�	�Ё-M��lE�	l6�q�>
�@bJ�(�$�1���,X��/s����?��A��B$�^��~z� ���!��݄��P�b�,.~�����o���MFL�H|S�:�H�a&갱��ʻo���8n<f�r��ƈ��.�t�M;!�s���׿ˡO�0�ǎPx�����&�� q��)�S�����=Lvd�~��w��;ϼNp����Rln�&17f��c���_D�_f���jW��x��!���u�W�Л�$�AU��b�+�����W��s���z�sg^a��w�J�o=^*F�Pj��f:��(ܸd1�H�#*����JT@�
�]w��ٚ�����*�¡C�ų�t�<���h{;���5�.tI
БF��=JzT��E��db��,X���l��� %5Ӣ��j���Y��g<��w� ����/���.7˲���N��{�n�}B
�6R(I�Mt�^��j���0�^/'��4��ҕ���.0?3��SN�}eY���P���eF�i�75�{��q1�16�t��ʪ��Z��1����@�t!`����W���p:�7N��c�r�����H4������c��f�X_]��Y��c��7}c�-J������$FQcQ�r>���$���y����vi��W�����&.����PUa��q#D8�B���˥$5�UH(r.�m��8J0�"��v&�ؽ'�#��1�ɘ8���{!A+��xLcj�,cfv6�o�eQRV�nȃ��Y���K�eTUō�7����O}��Լ�ګ|���x���ٿ�������?����g�}������`i�>Ο?O�场�N=L��p��177�[���h����70���RF@�#d$)�"�1j�fM�����T��ꬣ�,Cx��p�`0O�h�Xr��e�y���ܧ>ز���tD��1����9W���N��:>�Ii�xK�4�Dĭ��@���N�e:-Id�C���MYr��9�d�P
�*D����&7SՈrJ�LB5���^[F�m��W�'r�9��0�ηP^0��!>��(�p�	�D��+�-Q�"�oK.}�8����q���C�9$�y�Y��Ƴu�
k�|��'�7{SO�WopW>�!ߠ�fbU$�:���g��ދ�ݷ�$�a�E��E'M�f���Ux��C"Y8v �I�x���9�$s�Q�F8���D����&�ϽL������'i���W(���YNa<!�1�b�p_W�"fP���_���IzO>�C_�<Wߺ��jZ2��XSy�I$d
�g����Q�Te�d��x}���#ꊸ��YM�V���~���'8s�G!E��eC�iU������){��X�`�0�k��M&�JR*� �B>x�%�j��<ϻ����X�Y�x2evn�#G�0�N�NƬol��v��;�0M�6!a�U�5J�hfm�vm���#?t�J��,];IH��t��A�fe��nJ�CK������gXN���cρT�a��
uYR5�@��4a5g�y��sa%Q�Mp B�t��uL�b�ɔbZ�D1ܾq��W�p���p�
�Z���2�r��y��1����G�|�7fd��l���/����+bu���#U��!#tc������;҅��~n��X!�',�����4MM�fL�#��I�p�������"%q��E�q�qN�iAS����h��:�����\JA]W�U�Ԋ^�O�*�w�l��:�IӴ�i�����w�͞={(���d���
�9>���2�8�+����h���%O<�q~�g~�Sw�ǯ��_���_��gx��y��x���(���Ogn���������y������Q�K-Z)�r��!6���+�Sv����-!֊�xL�͐$
�,/��<��'�HFA�u�i�S���$ɨ�b<f��J�߁�U���uA�!�=~d8+�ڑ�+-��H�rDX���q]�4�)k���Ơhp�7t�b
��p�h�/k��`�Ԩ(&
c,V��A��Y�|���Mn��0�UzO=B���M��Or��x���d���.��MV��5WK֑��,J!:)P�M�#/�M�tu������k7i�]�P�1����,r
��9n���������|�-�K��i|1$�[�dYѝ�<7���<��2z��[���!�$�[�H���]$k������'�3�� ��tD�#�
Q�$R���
%� aI��j���osǁE�{s��}�TW메�ށ1k�x�~N=� L
(&�m�kkD�%���x�_e��Y�±w�^�HSm���>\eItaC�'\�p�HI�\�LY�kZK�� ��O���C�D*D} G)��u]�dYxvHE��'�v9p� {���p�����GC��癝�A	AQ�1��_��B�ڂ��I���	6Yk�0-I�sFG�4���������~}��$$4MŴ������J�y�$�73Cn��>�$�Ν��{�QW��Ȓ����C]7h)����.�Θf���\8��,�c|�0�j�U�t2�̻�p�����Z�]]��gtIz�zO+󄌣E���AZG�|t��TAB��G4���.S��^���ha��1i��)΋����T�?w����(AIE�&�E0T�X	��J��Z[��R�o�TP�zG�-M��c��$i�#t�7o�d4�f	�YJYag��~�O�"�����jU�Zk���w����a��53��6�yʉS�0����PV5/��2���|�s_�����������������������z�7�}��nr��%��HҔ��d}m���-t�PU%K��ܸ~S�ĭ�$�����5�l��#�TU�������1�ɔ�;����lm�����`v%#tҥ7���n�t���=�k6n�����?�M5�r�LG$�F	�0IC�"tU���k�iP۷�P{��V_�� �x,��$��k�A���-QB"�_c�?�&&I�Hhj����da��]�:��xa���Ho�͐�mh��|�ܺ�&�����}t�f�"E�1���ڰ}�2+�f��,	˾H����ĜB(���Ziʢ��%��-6^x�A/�|��k+��AM�YE,.����Fg?`�����r��o�]�J�.Q^�t�9�O6��,�����1S�h�yO�`�ƪ
�'��u��+Ϡo�"Z_��=�`UKģ-��Q��F2砩A6�?�8"�5�g�s���aan?���2��4~j��,-����I�!�p �Zr��((Z�4A��hM�{N��fS��9:���D���+/����*JH&E�] ��*L�i@��z`�ց-��iL�+~�V%eY�$J2�8!�S����lm�"S�,��QR����b�'dY��a"��)޻��S�<����C��qxVi��I��4�h_��ĺ���2:MN]���#�x�A�\�������--�g9��9�4����ɲk��4���$D>�)l;Im;�mBGc��&��m�'��$'7�2�����RL'�f�΢��t����<��%��5��RL'呹4>�w��xL��>:؏TAG\'��Z�}uY�k����m��:8!�;"װ�z��gާ,
�
c�(
��R�-e@7�U��B���]�JBP:�8k��T�`�,O9r�8q�2����ϖ��}�z�7�ts��4�=9��bsF � 	R"L��R������\���*�	�r�,���R�"	��v�� ��.������3��o:��o|�x��v/�PI�N�{j�{�=�{����wX.�*�M�ь�#._��`0�ijL[M��8��FK�r�b>��Z����붙2�<e���� G��t��5��qppĹ��9>��/~�����>�������/�������w�[>�����W���AL`B��y�/r��]ںbZWTu��ge��	Rog����DQ��s$���sH!��a�3;=᝷��'>�q��"�8!)ۖ�`H�NpMɝ7^c�HF�C�y�e�~V��P�gم,�{��_~@em� 8��d���8%��SL�+�i�XD�11)���X�{i���%<FxR\�h�R�z��Rz��ȃe;hҺ�<Xa��{ߒ�mC�2T%�4�Ōԭ�J`CzM�h-h�H�y� �HC*M�.HdՊ��ʯp�[�bce�n��p�O�'�v�aO���ܣ��<�{�o��Ĺ�-6B`\/I�Ez���K"r�ٔ�>���wh�g7(&�7%�� }TKS�FuћͨZ0���������1�*��H-JX޻��o����z��Ђ~���ʳtK�!�!���e���2FRC[!| ɖ1,o���/�Su��GZOp�V:*��Ž�!BKT^���I���Ҷ��C���:�}�m\gQ2�9������8�RH�p	JF�{��q�~�����!ڝ&`Ҍ'�|���M�9I����M��x���\�|�[�nE
��C�����n(˒�l�b����u>�g�B�3,��$I)����^��Xڶ�iJ�ajPz���O<��]��^{���y��d��y�ͭ-�x��}�m�����$+�;�q�v�)���)c��������R�GC��}H'MS��>���8wa�FuFtB���/
t������O��~��Ά�� �����	������1�;�%��MUa�8�������E��^��89>��;�2��|_a���D����:.D�T����߄��Bb���|Fc=B���Na&�ҔAZB����L&c&�1'''{{����$I���	7o����{S����n�L:��OQZ�)Y�1���ܡ�w����tF��|�K_䭷���x����/�6��?��L����pp�>{{�^�������o>@(I��x�b1��5R��?��D����s�Ċޣk��6�Y�!B��(����o��#�����d+��	��˗9y�6&$Ҳ!4[2���8��R ���A@p���&�K�4�4� #�iq¡M�PKT�ZYJ'��ce<�-��+p�8�ֲ�f��m Yo1Q�]��r:r��`u���!R��
�	�R0�&�8�$t> ��:D�p�!�	�$��@zp��q-��sـ=�`q>�$������I
S�
9 �X�g)fG��DЮj���B%�z&MC�z�1�A����d��^
��aTK*������K�]�`=������d:EF�ϸ	tZH�e�j`��H|"��wQ25����ԧ��$�+=('0.ޫV�� *%�w�)3آmq���=�����D����!�'S�Vxb�B)|��;K �DǤ?Z	k����R��I��Z۶�!IV����t�3�l��}���)���,+�ԧ>�O|�'x�?���Xk9wn��x�s.V⫒��(���pUU���ψX��4�'��hI���YA1 D��X.OY,gx�Ɠ	�u<��\�������S���ܹs$Y�'>�9�����u;t&ɨ�U�Q���aj��C���<:�ITo�5�Aе��ii����_�#�xt��4͐��&�6���DJ����YBn;�m˺y?\�ȑ�;t2<����"��@�ۀ�H�B�xgyp�.�''�IB`]4�B�j/Dõ���X��$z�1�=��	�4-�@׃�\�ʵ돓f9wn�F+�h<�i�]����&$I�x2�lln2�Ϲ{������ޡ��h�ZUX���DJ-{��`0`8!;�Ԟ�邽�=b�x2���[ܻw�4������;o����	�㇯��?�!^����}�6��/ ������y�����j���#�A�IS|�i\>���k��9y�!��w�������4�k�'lm��9|p�zU�C���4G���(�~jě�{_�	��t��B@G�Ϲ'�z]ii�A*�'�2
��pJ`����h���i��E�=A�d&%���@P��$T'��� 2����!����a���E���2�h<A��Z* �c|�̕�I�d��5�N	v�0���kIg���u��w$xDYR(I!4#oiB���[4m�es�Q>����xFm;��L� �MC+��ޥї�Z���1놌� \$	��*T����ø
�Y�QD����6r�IA�����)$`�n]�,�֡�-R(�Ԣ�O�t`;R!�0Ȱ���2Z{�vl��@m[��X�Qղ�Z��=�/F��}���#�ڌ�B�	ϝw9>>B���!x��3�ժ��BB~Z�,���jm�����>���dz�h��x� ������b<������M^|�~���7��W^agw'�;h���.UU���s��]NOg���XSż��+M�PW5f��d	�p�p�A����</���h@�LX-�4m�tz�r�dw{��x�xCQ�|�;��ƭ[�����>�!�ܹͫ���֔�S�!�5��ƑD��Ɯ!�Co��n�	ה�2n� �x��H���7oR��L�-@`��ن�3B�Q�G�Z�9�mg�hx���"@��?�_�����?�T��^�T�\�{!�{ve�T�3���9M�CĨ{�%�ߥ��d���A��uxo�Z/^�69Xە����"*�H�ll��c>��X.Y�V4UE�g�_�����TU����].]���Ƅ�(X,ܽw��9�h����
[WQ��Z�
Q���,��8��UlW��c.]y!���O����+���1�`ۖ��ۿ�%&������g�{��W��[������Ň>�1n߹�|6�jV$Y�i�m�!
fx8�ԓ$Z�ڦ��������-6�.C�ؒ4�FI�w��ru 6� �!�N�����݆D�H�&����+�R����>zv��y������#��4�RP75�r���H��:��@�
�~���E@�!#XND�Q��U`%��-�Xt"c����M���IN�~�}-�pI�gv�����u�R�k��Y� �՜�$$�wh��x{�����Y�¤��k�\�0OP�����[O�M�/������E��	��������4!�ID;w���> �Ba^@��GH�P/4�DA���HZ����u��C��F�b��[h;|�D*�T��{�9�b���"m�A�]�LeA%t:��H� ���V�x��.���X�ŞV��W�2v{����� k}�ȓ$���G?ʇ>�Q\�x�U�����>�A�Ihz��˗/3��J��1��𐣣c�!1)�"���D+svf��k�u����nS:���7O���ޠ(2�ߢ��4MIVd��̘�'H�8><"�<��Sܸy��i(���ß�'�w�&h�`8�نr�<+��R}p7gV��J#K��#)%Qڂ�kGiE�%x�9��;�n0��:�䵶�h�јb<�L�d���fC�=��������)�]�����>�F�)~{DQ����$�@Y�ȒD̞�6�v'Z�z���͡gq� U"ZX���q�X�-����&U��s��p��E������pȓO>I�$<xp�<Ϲr�
��N����� dyN��8��*.ئ�\=��|l����<�w�f/^��^��B������������-���p��ڶ�����o�_����$ܻs�kO<��g���K�/��O9=>�\�p�������!��\�h�	]Α���|�G�T�!���p�k AK�x<၀:X�$��al@X�
"�DD�/�}�X%�C�p(�KP�:��Ȁ����g>���w��H`3b�fpn�����`�n�b~x�0H  |0�����,^;��H�F�]�� ^t��N@�N#�N��Ē�+�Q�F���3$O�@s��Aה(_B�('�\�
�
���������%��v�4��'>��?O�5���%n��*�Υ� UZt�ǹ�u(��j��QG@��h�2 �@z	^ ���Q�b-������u����:�c)c���h,�B!�H��(�>R�Ђ�Jl�(Fh|�"md��Ϫ����Ǻ�]���WT���i��KWX�H����<). ��-�L�ݧkZ��;�I{۝%�I[�V����W�>&I��s��:5�rŀ,�onq��%&�Ng3��)�����&������k���١�*������߿��*�����ZD��]�G/�kjH��^��C.\������ϳ����b�O��O��,9$1�wz:#�[�Ο��7��Vdy������{�E�y�m���02�D�B_���������^�6�)4�u����^u�����;������Pڠ}�r���&>/Ȍ�UJ4�mive��ж^X�H�����3S��!xUfR�d��8D�]�r:��y�F�-$Z;�����˾^|��9��]�;���(�"�{��O=χ?�1q^�HE9�s~���]V���dc���{�m��\`gg���x�ͷ"U�E�� /�mG[�H!�LM�(/����`Rƣ	Y�#����KH	xG>����d����'��_�Lg3�d�o��o���$������l�RG�������W���dDjDԙ��>���x��S:�!��4��9�R��G��Z�隚��qt�R
]�l����ۆ�k��C���"*C��ӆ@&��M_�!���(�%=ʃ�Z�"1\��G���L>���1w��u|k0�!������<�'_������2�u/�S�.��	�O�@�b�Y�z�+5V
,��`	�"]��
���MS*��T��B?�8�C/Pw(MBӴh� �����Xy*#QZ�v��u�9�भx��K������!y��k�������Wf/�����u�D��D�j�i�Zt.�F�8��=�� P"��� �KpBR�&Qx�)j�r>V�֣����4Nb(���'8�HB�PHaA<�EZ�l=;���]�>�h�"BF�sC�,�ZX	�s�8\.�6"{�zB�!���(g�o�۶�Dc[Uڄ|8��
!l6�G���T�5�s0�ӌ�l��m>��Op��'�ڐ�9I��Ci�_�O=���	W�^�kB]����9�[L��xp��{w�2_���!ph��"�%�y� #%E��ey��v6�y����_�H1(p�E�wα��E�cB�����M>3٠�����pB��fw�<W�x�;7�ÕK�V��'<Z%�'��H��&~�fEEs���(Гe��h;K�6J�Z���aT�Q�IɈ��GcV�A&��/��VR\�ok[�c��[��Q@���	I(���
�
��v.aE�Q!��@P������}@��H�P�dxkize� �^Dt�@�B�R<J8��,M�"EA�Fd�&���ϒ�clW�5q���x��<�I�q:_�s�"O<��p��=u�ɇ��x�jYsnw��t����.8��BT�J3�4e�ɳ4R=|l�(����A��sj�N��+ן�ʵ'x�C��u����;o��o~�K�����ԝ�����s{8�H�\���s�9zp�TI�7�h�c6��Z�Q�\g�Zb�@	MU�XU���!27tޓ�`�A9��x�y}���q9J�.R�<���r���U	:O(W��`ɴA8O�E�@'bX9I�%B�Ft���aG#��]�}.n\�ucN����p�ß#�ɟ&\ ��bF4NS{I��|Lm��$aS%��S*�)-~�A�Ȕ����1�8|j��Fu��R!(�$�	�c6AB�Ѯ$dP���ih���,�	~8�+q͒kÂ�|@h,U����u�}�:����9�Y����7�	�R�3N6���j錧v� �B8<ì��|�R�@c��a��F
 C@��i
i��V��,��fs��]r\���eM�[�iñ����	��,g�F�� ��?R����l�����9�/{6��yu�!T/���	��-��=�X)�Ɉ���Ԅ�@�G,O�\}�"��v	���4���P��MM�E`��qF�DL��w4U�V�,�QR\<O�HO �ƐT�������6���iAմTu�2)O=}���מ|�d��wl�?�d2�ܥKTeɪZQ�탻#PF�U��t���uZQd9���$I!�y�F��I�d���#���4[;ѡ�\����N6��a����C�{�=�]�������8w�
���������w(668�Ͱ�#OR��Խ�e��_F Mrf���*/H�Bk��e�68D��X�{��!ˇ� DТ�
���9��V���˂`�w-�.��ż��
FևT"�:!�G(�� �xDD�1;9���R��j��h�v[W�u=�%�Ԝ���Z�#D�>��$�nnweR�r�j��*K��vvwXU'����j�Z�L6��6H���w�(r�4��k\א�8O/ҌAV�ʼ�xi:p�D�˪�*+�u|���1�I��k�t�
W.]���(_��/�կ}�͝]^��OP�5���x�2�L���UܹAնhc�IAP���Cz����{Fo���UU�GX�(���mT��/��m[��eY^P�f� l�A�I'N�ú:�COg�h$2(��j�o]��]��������7�[��x�g>C���Mi�S�;��J���a���є���G��~�'y��g9��r���	۟���|u�:����or���E8<f5=E=�8��>�+F�Hl�{�.o�&X��2�<�S��T�g)!)x��Mv��_�'~�s�����|����
��$Y���KN ǻv�@�/�̙�����/W���q��װՌfP .�����ؓ)����᭻h��u�qv?�je���+�X�z���_���.��c��;{���g�{�q����w�o�gX[V"���0�?ù�~��l���7�����g%�T�"�x����(5J
�eG���X[�:E"�x��.�U�r�6�ם�p�������sm�͖��F��m�N���D�΄�W+NN�x�It�Q�q��4)�u�܈��Fg�uU�d�0���lc{��(���akw'���0��`8�����o�EY7q\$$I���9;;�L&�^���ƛ���i���Dc�������1�(���$h�������@4+��4�Ő��X�Ts��u66�h���d#����g-*I����Z���4���dd됩���$:k1RF�)����7��	t�rzz�|:%�Q�Q��t�p��)��D�H)�� ޯ�s����(��~v��rȤ��$!�r�1Q��W]������Ql{8W��+�����jA�6�a�Z0%r��C<8��C(�`R0����g��(
Do��4I�rn���{�{E�w������.^��r6e1=d1�Z��Β&��$��`�Di1k���ڦ���*�4ːBE
^h��m�kk�<��g�a8���MS�lmm�)��Y�Q��K�=Ʒ�ah��%Mgv��%Rk|�4z����l���/��`@�E����؀3��"/�KI�O�~�F����#DT��x	]�c�"�
�h1B��Ђ�������B�o�>w������k8|�����?���;~�%��P<�|�s���.ۏ_e���'����:%5	��&����+w���%�_�i�1Ɂ����r�_��,�F�et�1�i�%��.��������y�|\���ǟaot����W`�`��A{oEyoNq�:/]�o����᫯�޼������	��l<�?�)��0�n�[��,�w��k���<�� ��s�����ps°��*W���7뷨��G#�l�����>C3I�Ҫ����礲a�����_�|�9��a$�էO=�K�ͯ
ť>����/0����	�>���]��>k4���,kʘ��L`=C�C��T/y
]�2��@$	I���Qw\C��e�X�g8R-VTU	=��[�N�Yb�}����۶_�Zk�,�
q!�^�!�`����M&4�E���خc>�1{��i�p8d2��e񹤈ΆE������d���o�1$Z���޺���IB� %�����c����rJF�)��%`�X`��;OQlnms��4u��<��&M�llra�&t�6�1;9����$dYyDL�#�.J�f��<�!�;�4I0�����"�ѝ�����+Ʋ�iӟIJ[����]���
��!0�DJ)�I�iR����GCD����"�$+2ʺ��-�~.�5�)nJ�^� ���D� �:���bPp��u��1���j���>���$�C�,��Tg���ۮ�uZ�֌��Pd)E��hu�|NC۶,%�SduC�v4��k{����X��I��d-[�|�3���;Ν?ύ�nEm�`�J����`�j1'Ҋ�|e׶�!J?��$w��g#���i��\���N�1��RW1��>:����|o>�>$!�{�PF��������V����8�(����{�,R�}���I?g<�AZ0]���_��]�hJ��4:�S�l�(
f����p��U�r�bq����jC����ӟ���xs��e�٬s��!�Əw���r^rZ�|������"8��!]à�?�"������e�3H�(��;��O�皆ᇞ繧��g���Nw/r�׿��[F�$���e�8�wo@�y�ɧȞ� ��78}�>{"�lDȇ �ɒ|{���^��r��/�C�}��?���a5=$����}^�����<��\����5�h���1�*��[l}槰_�����m��H�Jx0��9�vtMR�v�^b��8C��{x���3���r�Z����F#�����_#ŗˈ1J���A��n��G�C x�V�:�2��u]ۃ�b�+�3���9��!{��!�<�\���dB۶�?�ϥK�{�)Y�N��V��pHf��`��)�,�w����h�#�n���Qٲ^�8==�,WQ�a�����0y!��ьJF��r��{w������KZ4}��K�.��2]�PZ���{�Z�Tq����v�E�ҸR�31�5=VI�%u]sz:�Ł^�"~�@��)	��.��e	����x���iE��iD����J���c��*�Τ��-�u�ތ������mR	>{�QR�$1
%5�ɘ��-�"'�3t����z���B L��lܔ=N �6>���k(���xL�Z����{$&ڸz�!Rۄ ��)���n�:ۋN�d(�����J�Z׋�8N��<���+ʲ�7o*��ePlmos��-�u�i���z-�JD�g-���$I������a����n*�.j�/V+���M��2�k�M-֝�N@wQ�FyH'P>���9N��W���x��{�����'�D,K�|�C�Lr.����-�K@4Rs2`.\�DҤ�J:�����4�a4V@�%.Q\����������ʟ���w������{�nθ��O2 �J���}2�3�'ټv5Ί��,�-	b���9B&����|�p�����Y���[���+�{�*W/?��O������j���pB�$��>9)I�J3'H���}�[|��~�s��9�x��y�֑����1Nwt���ÐS5D�c��EB:��������<�{�����@~���O�ǿ�����C�,x�w���/~���G��f�4�iΒf|T��k��Έ>��Y�:�D�r�b����=����&B�^^�s�V+NOOH1�FC��Iz�4�*kr~�6�(б��J�Z�$Y>i�<�s��x���xߓ�X,���X,��١�s�f.��E���S��r6�$JsR�$J3��fsd���Ͻ��݉FJ<Bkd��ڎ�|�rƜ)?:�b�y�1IQ*��,���<8�_����g��@�h���y^N{�$�.b�h�i��g�����M��I}�e��R;G�>��:�b���ǂ(\T,Vx�	�*�����g�ݿ���'�ú*T.�Bj�C0Z�;؟emB��`�\\ԝ�4m���-����J��u�ij�JX���c���)��z˃ш��٠��4]L�4%ˋH��[Gy)+k7¹(-�%i���[�dp4Պ��4"\���Ժ�Z�(�P�B�Q��;����օ�,�x�h�������k�C�� ���cNg��m�`��U�`����+������sz��3;h��{L���1���c��=uאH��R �q���%�T8k	���(M)�גb�m�c�`��)A� �"�Sx��L��qTG������]f�u~�~x��~���/q�s -H�E�VP54����(rkL��>~ P�)�nN�:��^b�k�'�F+ùg��|�q���?%=���%j�����;8�1X�H��i2[a�#gl_��ͷ�"SD���iVP�{@yx��H8�Ɵ����-�	�rE��؍�᳗��'>�]�k��!/���Oo�%�<�r��C����#�jP��4��v�����]Ҧ���,ؖ��ۼ��oa��S0�K�e��7_g��_�����~�5b��繒�����T�
�8�S�fK��A+E�^dH��,4bU��p��+��T����Z�LbP�s���m�X�G�@D��ZC�A���<m���xa�V��K�3wF�&,J��,�;��AϏ��"�i�=K(�4g8��2�!D�A1�{�Ng����b4a�a8bt���" xU(��Dő������0"\�I)�&�Z��"[�4u��TUEV}�,~�q2�2@ĳ�E�����7op��-�,!�S����5��4�6��4�8#�:���j�D�z)�}�u-BEA"4H�����k�y!.xdjH�Տ���(�t߻{߈Ž�z�R�{%}1��\����n�G�i����TMCg;�� D���<MI��D�Eed��R���#P5F��,���![�q�Gl��M��
���6�-eYl]ٵ��Z��D��8��,ʪ<����"u�#��մ-uےh�%�,EǶ��Xk�>�����
� ��8F�׵�FCꪢ\�ؘ�"F)t�1�l����l:�\F9�,M��u�v1���FJ�2eHAӶx M�r���������j��o�����#���'d)D�K�b�q7�|���λ��DL��x��$#�-�+�;7�Kl]�����/B�i72\�0�H#�}�1��&3,E9g4���T��13}�&� �g������ϑ��^��?�Mfn�(,	�b�=�3?�)�_�^�ï��~��|��r���{�,K�U�;�ߠ���h���fk�I�3t�.]�g>��=�"׫{L.���+��)���{/}��W�й��[o�L+�z�"��c�UI�eX#��,v�b�.;��fTR�y�[�\%�0�N0!e��A^���pt�6�o����s��'����eo�2�քp<e�oSb�B�"M	�$U��N��j��Hm6
@�D�?�:p���b]C���o�K)���Fc������tm�K.k���)�3�C���V)�q�#��봟�M�%��"��"Z��~�:gAD��|���������S
�Z���CD�����`���E�&R!��!]����P}�/BD�_���`�Qu-��컐�<Z��!"Ҵ6X0I4X��qno�����.D�;����Ĺ���[����A@�t1���q��B ���#8G��ύf�,;���l�GƄ�G&etLF��&E�*���}�#����m[������meD?���i�↖��t�`8 њr1�[Zq~�Ά	�_�1Qh�d�"�fY�(�^I.�oڦA
I�$1{����HR��M��bQ�.Z��y��tJ�Z�M���cWAI,�������5��<�C���똷n���,
a=JJ���.^ass#�!�Y��gv���=� DTo�%������B#�ǑD�����	!�g-P�g{k���i4��yQP�lg988�*K~-k��[��i��RDD��
�#��ip*`�C8KX�r��{��{�V�G��*:��<F��������/�?�����*��t�M/H�����>�!�=O��a6C,WU������W�!ŕ}����{nH{�߽Mz�m�7ϡt�ŭ	O�?�����kƗ�2�r����_"Q��������e�N1b��Y;\7���+��1�g��&!���)_�*�o��u̿�u��<�$��Ǥ�."��5ܕ��K���Z�K)\`G���a� K˨�ا?��0!��TV3��7Q�S���o��{dy��/>��
ڗ_�}�M�T �[@+IE��M��m+�T mK�i��5�d�:�1�ݺ �Z��k�4y�$�W+\�`�,bc���w�hQ=b<�,��X��*�s� OS��tM��MC��$�yD��TJ��q?��Hy�yV�\.X.�@�����y��}ضE�FtuC����y�.�i�DKٟ��뢮@��!����u��C�Qs	0�@�]�u?
�s����W���`8��w���"Ǉ��>"ڵ���g�����	�V�TȨ��zQE�w��h6�Ӄ�b�����!���I�����z�t .N�!�|p�E0V�q�(�(T�u�����4��b��Xi�zPK��5�=��@�f*&�Z�EAZ�^bt���pm�:Cn�X�
�p�s���p�h4�vF��1eU�XK����$	i���]Gݶ�bL.f���u�|��ԡ�l�Fk�<C�X��딛eڮ��z�ÞmpH�(|@h��.V! ��	Eӵ��C"O��"c�Ū����,qޓ���F}L�"���]ڃ�D7.�t��DG&A~�_!o�br�6�.�-M��}�=f��˨������;�8��/2z�]�LY�N�y�Q	����Ҭ�~��PǷ�x�#���q�×���k_e{>�H���oq��G��\�|���{��1/��2�O�m�^~�u�c�	���핥��#�����7���1�yA�Z���x��+��$���7FL8}�U�|��X�(�&����o>���&��*�{���S,�7��E�0��&Ϟ���~2E}�-6�"W�����'?L��u�[��x���G$w�sYVo���o~��C������!w~��<�r5׬�~���ߢ���7�k-��`Iim������c�uED���?�X6MC��19a���F�Mϒ�\�5��G� �Q*�FY���w1�y���<�I�h��ǌ��?/@):�0ID�K��������g���B����ߧ�:�����|8�}��� �-��4��"?��xd?����^�yL�����pz:Eq|&��7�B0��s�&R*���H�HK�Q��9\��g�s���(�
ۖtu�VI_��{B�v�m��c=���#i���@��>
I)�R:xA?�9�0�쯬۶RG�Rdy��Α���r��5��
��Y�P�5i��򇝃��H�X����Bir6���٫��3hd��G�1.]�,K������"��W��T+
�#��t5���
�"%M������B������b��(�V�<ˣ�Zb7�Co�Zqx��R��Lk��]#S�v��paR����+-��F:�飯%������.+���s���-�,CUm���LOA���Q�5�<���]:@`������u�Hq�)��>W߹���#]���EJp��W�����m,BIג�Ӄ��֛�y��}��!�0����!�ޑt-�j�b>��߂\�a���$�,��bu�6o��A;/��3��緷����_�}nMO�1�.2vRó;cv�"l��
�=���,����H:Haq
�){u�f��	订�ӯS}�{xm^и�.9�����ݘq��y��Iv��sMB�����o�k�݂"a�t��W9���	�!J(���c�
dװ�z�_�&�_z��뭍��H�"H��7��/�춆��X�!M�E<�����l��n���m�5�lȲЭui�}~}N�pD�jb4Z+���=]dlzfF۶�4��?kTo�,���Nc�O}՘&)�n�^7^�%ʏ�?�M=��i���s�$䃂jU��|k�GnJ�MB�+�����2�#/���]�=�-��$(���x�������:���;mG�e4mK�wR# jՋ�x$�l�{%�:K~��O�:G@b��󎲫Q�GʯG�>�k�=�-��_��SJ�N&�'�l��p�:賵GОȊ�����I)\�x�:��3�Y$�H" F�FRI��H�����:c�Hܘ��=@D������F�!.@Y�����bC4�> �CY�n;��t�a���k��e0����!�R�6�/�9�H�|�4��P^,kZ]�vx�ɲ�#f�{��$h��(u!P:z@�~s��:G���ZD�R�V�q cYemG]�x������ 8�|���!��]�S�V!�T�%��DI������C�5uM��cK	�6��$K5�n ׈�D�+hK�f@�����G��th0�S7��RK��W	-�ZF��\X��*H��m1цU7g�8E�+��\2Ƴ��C�[RQ�h>Dp�a�����y�Dܾ�X�t�E�����,aTw��.J�z�/<�\2l=�Wd"�i[�ƀ$$ �)��$I�r��4�~���%��`�(�,���Hl�XԄ�S	��@H��[.(�IfH���U��;T6�����OIH+��X���8���Q�ߛR��������h���A��#��,���"(I�:���Oܗ�k{JY��u�i����i�Fs��y�c]�h��|��Uѱp� �i��Qߴ|�!#$<�������F��/˒�;��s=GW�A�Y�ȥ��>�!C�ѫ���6ʻ�������ϦEt�{���cZ��L&�<�b�JS\��|8�?.�j�h��e�="(|^�W��"ơ�d.{��'H�Q�]�(]��	��$���z��Cx��ǀ�\<p���>�=]U˺�m[lo"�$F���D�tO�Ӛ@D{:ۜe��2L��R��9�Ra�mb5��t:c�v��ʲ��ƌ;"��,'A�f�B�P��=4^u�󠴊��y��)�A��ք��	&�gw+��8�b��;�&�OeY�;B���{s��ͮ놺i��C���,�g�2kmoiq��1��G��uQB4�$���K%����HSV�Y��*�ϧ��� E��!�w�@���N�i�Its���H��0��4t�Cd)J8D���t��WP9Z!Kh
�L�Β��L�	.u����Y�-y��u��t��>V]G����6�2TՊ�^�UKr��MB��iZ��aQ ����F�iA�'u�R,��k��
�┐AekjH��8A�A�$r�۾R�`4"Mh�f��N����>!8��#����5�6K�I��.Ŗ5�ʢs��ZtH�	�a�d�Zc���B�D��:6M��|4��Td�h�ǚ!��N�B�#gď̄]�2�P�V}�Y��!bҸZ���
g�L�;GP���3m�Z�1!��"H�~�+l�}�!�X,����HC�ޣ��Ҭ�T����M�h��3��������jE�:l�F�W�}�5�����C��:1�������X�>ʲ�v�`\��TU�|>���˱�� �� ���ܿs��p�b5���"$���a��$	J�؂w+�9���|��ř���\��G}�UD��j�:��	m"��oѿO���+��9Q����t�o������*t�h��6n4��Fu�$$J�6��g� J���D�U��]K�6�<�e�ZQ�+l�"e9���e�xsBdZf�[�i��֞�X���M�	�L�����)���zOfB<��,��dY�xc�$��5a4�$B>�>��<��FA|l�$�!x��:��q�Fμ�nL�gp��E��1�1=������P=���v�c�.xI�����}��xڮ�r����:ъ`7�\�7y�y��.[V;Lp�x?�TT���3(R&`=Y�H�hl!��-ao{�A��=Zh��&����e�'�$�;�a�W���"6��DM�m��*Q]�}�M���_ĴF�i�Hh�t��М.��9"X24N$,��͇�<s��O����K����4�0���#�%�����L
�H x�LdL���v�C�	^�#�VJ��e��Ks�
�?�)�^|�=������׿�ݯ�1��-���j��!�����
G�"3�t�	�a�C8Gct4�TBh[� ø@&$������-]׏��3�G��JJ���^.�$i�ZEmٯ�w���Y�Jto$%X�Fs���g�>��ܺnٯ��<G)E�Ԙb@��u"O�^�i���y��S�:��&'g�QD3��x����`���Q�����;�A����½��`8`s{��dһ���}����i�����b׵}��)�*>���&MUQUU�Z�q�ñZ��I��{Q����]?Ԡ"5�x8,QT_�y�ƢG9m�PU+k�m㊏���r�ozܨ� pB����l��*B]E���
���:��PZ��ߖH���
���֖a��|@*�h4b��l� ���JBB�:lk�;ڪ��!�ބ��4!HAY��!M"Mm1_0M�R��m)�KbҢ��V+����ਔ��#�ʑ�lnlF�j��z���Fl{')JF5��$B>:D��@��^P>8ڦ���R�}���$��JV�H1˴��
�s�p��M�������D�j��Ρ�68К����I
��6��#<�eUQ�-c!c��{-�~|}�@���^��B�x�	D/8$*��'H����h�bc��!H�q�Б��$.���)h�e�%K�q��	��	�MB+b��Z�B�S��+j�o~�����j�MG�F@�U��m#���
��mK�!;��ӿ�>�q�R�A�	Q�)�1-BV���7^Ev0jZriH*�wZ��0�#�EK��"�aj������_��O~���%�`BhB&LFW�<C�싼��������ۧ���aD?� a"8�֣4"x0:� Aؘ����'nA�X?�	�}��"VD��C�=����R�E���j��6x�6��L^`�%_3|�I�w�����/�{��z�z�7��ap	=}Nңܣ	�����D"�C�5��S7&�Q�M�Ⱦ�Ah:ѨD#��kAUŤ�*	���y�2Q"�(�Y�`<fsk���1I�	>�U�$ygi�����*�P�"�-���^�"��Q�K��O�NOiێ�nI�$�Ȟ	D܁�s|��� z��!:[z���YCU7��:�	A�S��mR U��l�I�I*�h���#(���z�t�k��  |e�~5�.	:!H�*R���bT E�%[�Bf�!��l�A�oQ":�!�ilI���!z�KEW����+��2���$�)��1��b2��6-MUc��o��J�׃<�����s��}�i�czT�o^"�AJC��ii�cYU�c�|@<D��Ŋ$�@8�� <�jA]W��@JX��y��^��<w�2��9ӖK��b<gnt�E�@�#���,�w��c�7��x�V8$�UI6��i<���mW�ՂBʲ�u��WZ�*Z���2H�ēx��
��*e.���3W ��$P�C�Z	��֡�d�Ax�����F/��<M1�v�����2�&'�5Ȣ@��U1d�*g"5�"�>.�����C��=��L!�����m�3�*�8ᑾ#�<��� ���X�V�`�	TSGUD9�A���"��KG��`���>����,<��Sd�Fx%��Dl��y����|Ƀ�nS�l�µ-"(�JPB!|�5s.Ҝ��v�nx�k�sD�KA]� :� �s}�P=	ܯ�"V�q�}�	��'M�vԫ�ł�`D��()K�ln��C�	�+GJ}:�:�6Φ�����X,�F����m�G#�s�NO	�Š%b@OҘ���ib�#���m8>9F ��L��[E�T!(�H��s�ѐ�m��fg���=���!��ѽ��ѱ.���>���J�[��9R�� Sk[������x�ի��(AJ���T4�傓�V���"R�he�: I���i�"A���H@��A�!��j���eS��F��3RR����TY�F�<:Y��uqFK|?\變��e:�R�Z.��
�b�F�>=�#�b�1AHI�jpD��X����UV�뺗�$�`���,��FQz��#���-�)#�\������/q��E6�v9>:d{k�$���,K{lԍ7�0�hQ)M����^���J���u\ܓ��Q>�6->�e���i;}\.�s��V�����r��u�;�<������4I)gS֪m�V��'Iz���$�:+r�FF����4M�떲>fp��N����%Z(�д�e=t��b PR����dt�h�㉳I?�O����7��6}�3~������V��*D�� �eY�dD@YU�mG��RH���M>jjDבԊT(����Z *UN#�A��Cz�v>v��z�����S�Gp}Uk��FF�w�N�ޑ]�g���G]�
.V�g7#vI��������w�%�^�F-�� {�F�e{U�>�&��[/�*���|���g?��\9�B/!�ˮ_BDP���IQ���.��\,Y�f���N��f(E�c��t�%IY��8���K��C��詊�UT��&,W+F�(��t�ILjt�MB����IҸ_���9�Ŝ,KI�⬥�#�2��	�h�p<�,+��IR)���W����4�$%�R�,CʵNGL�sHe�bz|���}�:
�H�X-� Χ>�i67��N�<��D�@T�\{;�߂�x��h���7�QJ�v���Y��8�R����j����W�p�A�Y�N�{l]lw!xEhx�D(Cxt��[|��z���������U24u%���Qۡ} 8���xrD�" D#���`�vQ׸��(%{� I��?��_;��p6P��Y,W윿p���b��~��~�Ǯ\g�"��獎`R���",�dY
���_U�f�hS�:��ݏBR�!��7��L&����x�Q�J��6pzz�XU�4خ#MM��G��'S��������Z��pAE����m�@L��� m�M��Np�����)���e4�"Ρ�Zp��I�(gIPh!�"|M@[�(�P�s�>(=1�y����������5��(A�R*R!�� �B�@?� �R����R�%�r�+u��"C�)TBdLn���Ż.�;���H���΃�j��Z���8Ã�xg�A�]J��TB2y�*��'q6@�02C8��A���x�s6?�"�o|���o�
I�*�Z��$Q�?b*$^E��������k�V �����("������I���d�ەR`�B��j����]G����=��hM���w8Gf�$E�����zF4]��T��)�JE���ri�mŒ6�>x�`�(�RLO�lln���]��*�"?C��͝���;��LAH�14]ן�)�YKY��Ħ�{{��=��6J������b�h2f>[1�l���_������~��jIQ�NP� z��G>8���~��	y�b������1�"H�����O�}���������!�4�A�=��;�]���|Տ��NkY'"Ҍ�'���q����P�Tp��T��.��if3dۡ�����A"�s�~�vo��,H7]%I{���(���x���3IBF4p]�ض�)K�ܡ�Z��qn�R���'�`kk���{��|�[���Kخ#8���!�
��Ei�x<�ڵk����m�5�&"^��t]K��.�z�$�j�JFL���VEl�߱Z�899$�s��& h���rI1�6x�����;w�R��������Kb�N0�е�n����K`{��Q�	��H���{�.0o#E�m��,��cy2#���踤UԒ�H+D�0ht�?}��?Z�?\H�!~���w=����ElS:Zt����)Iti�`2ack�,ϱ.
�t]+S��j)����`4��$6H	��1�Zv�t��@g<eh���Z�����T�mwkoi���� �n4F\���U�h/��=u26%|TV��`��0a��i����{�>9�K[�����<\g���������c��q�5d���[��sC���DHG���F{�o���	����a*Hr�1��,I��4aPdg]��O�ٔ'��� &�@��AX��ܽ{ m����p6�;<<�k[���$	[�[��3�Y�4��G/���ol���	a�b���:����z�-��m��~H3]�f;˽۷8=9A
�^�����}��K/�ͪg���w��z�M�޽�b>�vk)�^�5����E����2�k��s���A�v4m�޹s\�|���]�����Ե-��ض�:9�VA(�֍��(�z)A����M@_;m�qR.�V�:e��)�mQ=2�C����8��)IS7,��(��/"!y�eUBt��	q��IB��h%�=�ҵ5]����3;99�	A`��$)��/��O|�������η��/}���Cf��ܺ�bv��mU�1ѽMG>l�g�Q�!���M߶��9�Z��5�[.������!���d��#�`�\��9��i?����X�4���LO��2&fös�׼<C;�h��m�Q�u�Q8�{f@]74mB��9A��0:� �ZG���L��[�''(���b�F�XMJ7��E-D��{!���x���=�� ��4�ƥ
���@��jgʃ�x�$T:-�F3�����]�r���^b���.GB��(�i������bI�<VE@�p��m�xo�ii�3� �@�Zʶf�T̖K���ł�bŬ\��*��ҡY*�� 1h�E=�8��?��
�A��^j����,����wZ�G&�/�ÚV�H�~�~�G��?�!�wׇċ�K���}@ͤ�[���S�Z�rI��G+l7�L�(�eIp-TO��h�{yh�V:z(ɏ�(Ą�9G[׸.v�D���Cn߸�m���D���m�������~��%�m�r����it���(e�(D��}�B��ُ�$]g�x����چ�����s����cn��.o����)��)7�{����LY�{�9�/\�����D^�ygm���)��<
ܸ(���)i���'$��@�v�;�4={��F��U� X�w�?`�Z1p]ޱ�O��Ůt�� A�Љ�r��uBtVI�z߄��O˽��AF�+U�;n���Z%~���E�ޑ���RiƓ�#�G���G�U�MV�R.J�Z�Z*��񐕂4M0}V��_Wܻ{���1;�%�4GO�5\��8?��X�|�����^�{��.��������stp�I5F��޽ͪ\�i��+��k9���<9:�[؜l��o}�Ǯ<F^D�L��X�c98�����,g:=e<ڠ��������X��ܻ}�"1�oZ|%%����8��+�o@:��C�H-qxVUEn4�Go�$ChCgi1B(lݱ�͑>PU%�b�H�J�A���4/�=> ��H�T=Dן����;��������w��O�ו��3䰀��F=Ny��}Q)�Z��tD�b���Q�"u�$y�2ʇ M��t�S
���8*82e��'��C�t��~��Ht��j+�rNZ����B��O�� ;G[6<Ђ��e($r0 ��GvKD��4Q:�F8��Z� ��x#�Y/z�	=�-�ޥ�-{1���Q�*}�.O�� �Z,D>26��,�.��n��qA!��P��s�'���єQ�OomDL��E�`0�2	�NHڦ%���pHS�Tm�]B�hp�Q��蔊�EUU�������k��2;>a{�h��@�FJX�?�[nݼA[����s|x��۷���b0���b�\�fL��O�vB"���}4�
�#�@�f(���Y�NmZ��8:<�-K���bN����m������NO����K��4e��;�Y.�&��)ɓ�AVеM�Q]/��s�'E i@��i����)+軜RkVU���1:����Ci���'���x����zQ"�
N��.�[^H�Tz��Žo������/��HP'e+�y}��Qz�Н����E�_"�s��sM�`���h4��W_��b@Ӵ�D�d	�u���0�S666������$ɠ��N�<��4]����I��Z^}�U�_�J1J���#5�4�Z���g����;��ӟ����7��_�5���o��/0�����)U����۴]�`��4��{���t]W�ޖu8�3�6u�bgg��x����bJ�Q�ڮ�4+�J�r�:7�y�d���1�0꺚��yp�.w�P�Q�'�qFصQ6S	��|���Ց�����6�Z�9G�fq�XVX��)ؘL�%x�`��D����,Y"2"�������)@*�J��Љxߍ�zzu��8��K=���� ��林B��F��"���X��`�Di���9|��T7E�vh��,Te��/��sT��)I��a>��҃ǡDD�+��MBҜ.�;�ʲx�]�w��1.(�����AEڏ].8���45�mȍDKM�9"�Z���Y�p�b4&Ã����~�v1���O��5��]�c��ƹ�r%]�(����e�F�2�<��� ��#	J�65I�F@T��X]_`� y��3'A H�J��QX%Њ@Y�� �P�����Mv�y����y�rԐH�3��=.]���������N�%��IH��Z��$4]Ďx�3`:����R�&x�i0�	�n��՗���?�Y��d�m�s���?��$Z��W_��j�����>���K6(@J����3?�R���\`m��OJ��&�ڶ����%Z���8����1㺎���㋪�D��L9o��]�0���G�Ng-o�����/r�����U�J�*W4UI�&��M�T�4����(���Aж��d���YVU�Ͻ��d�wBiÌb�sr�Y��Bªs�k}�^*﵎�U����&�C��S���N�'���M��fs���B����"*���˼���b��nj�Vg*ER���|F���tՋ��q�9dph���&���o��͛<�܋H�eη�����cW����$_��_�\.���>��O?�����s��=��/�T���a���&M�2=��-x}�K�$���@]�4M�ˤ:[s|r@U/0F�\��Iřy�is�SO=GY5Og<��S�������o���8����18G�W���?�[^W��E��[��}n���T�4�J�*k�_������Zѕ%���R.f,����ڀ���Ӵ����u� ���B�JM&�'vS��kn��	�R��`��n@X��� Ph�9�-3�� CB�ml}�����C���@u�W_�!�n��'�A� R[��1I��ה4H:!�
P�qQ��7��[�ɗ�%�x�V��l*��y�?���e0����j��b�ֶ8!p�6h�#�}��[j�;#T�ּw�_��7����<~�2?�7�:�b2B
�h�;ڶ�-c ̔Aij>���X��6`B��E�2������
�A�`9+��VB�!�`��a��f��2�B�B��!�rZ"˰6�����:�r-�8Y.������(���bQU��E(���E���(1����kd����q��e�����E���Eu����ǟz��������lir�a5�a�b8�y��7(W��k�q�滬ʒ�i9��rxp���	��o-"����$J�%)��enߺɗ������T%J��
o-w��!����L�Sx��"�6X-�|��_��w�EII�\b�f���#?�hCQ�M�]W:jޯ�]C��N	�Z���h;U�֚���`!E��7Ζt�SĪƮjʎ�G��2�7����*���W1�{�qMsL��M�<�V+ڃC��$L&8Б:x����-����DspxtVŭ�������Ѻ�p�&DUq6j8ۮ�u-��ܸq�+מDgy����T��<c5�#����+|�����o���~�ãc��L�cU���ˋ/~ ��tF�����,��3Q��Uc��H��%e9�UA����aA���U��ǟd2�d6_0�ؿx�׸�8�����k���AF�2@$��������h�y�*{:p�7�B���Q]CY״!]���Og[V�Sd��������tdJ������EC�8�Ou���!d����Z�7���Z�������3vց��)QY�ͪ�6�`$o|���x凸�#�ŒI#��mn�����H.n���P��<��g��p�?�F9������$M�H2u<���K�����]�i���/�onr��y��������S�ۡ<=��˞�'hmЩA��$���y:��h.4c�������W�ʿ��������SO��i��y��	J"���J)��	]9��#���U�N���Vl�U�d8�6�����Mvj���� �A��!��}�f�!jJ�MI&��s�''��F����lJ��	B�d��/`�>�'�9&ь'�ޥ����5�۶��h��0	�gAgmL����d��h���#����ٿ�����C������hx�5�gv�����$c�hMI<�|ע�-#��;�'���<Mb�q�/�	Teɭ[7���d4Q�+��0J1?�2_,���Un��.{���W^����l�;���믿���1Zk�U[&:�h�j���ڝ[Sݤ�-1����T�"b1�����!%W�_��:%����kf�S��� �Vs�[{!���e�y?\變�'(MH�X�k߫��SB�9<b0����B��M}l��0�N��t/l��Ѡ$UAl%G~� 5I?�����g�|AY/�M�'��i�^��.\����٧�x�⺖D+���mG����\}�I��_�k�������	�p��}<���K���\������JS�5�ł��#n߾��{���\Lπs�"��1�J�eLPf�S��)O>��_{���)�S�<�1�x���[���W���{���[ղwF����b�(�1��?AFjC]6�8�*�F7�{���w�V�c�jA ��Rh	2D�kX�[El�F�QD�*�"�X��}��r�<���3��Z�B�h��b%S�1�����{����d�\�y:���cd>�n��|�2��OD_jkI�!�2ReI�jY9��>��A�i� K4$� ��koP���ٿ��l>~v6�{�&3|�O�ť�w)v�h��4�QB�ei�����k=.(��6hL�!\�X�i�҄�?�O?�$O=y�;/����w�g��:�?�>�w�=.?�4�������q-����1ZAuZ�S뜃՜e]��"��&&4�C���@�%���x=�_�B����&���e�h��0I��,�6,�wo�$�p�����ȉ�GJ�ūWnl0�Ƕ?�EURV6F㞦��"�v˪B�g��y�p62[�����<?���<���`r.���R�����yp�>W�B��ܹu���	;[���֛(���"�	�(A�%x; K$�`��XqJd��g�o��}%����6��SV�9��dwoB�ޝۼ�֛�i��˗�$"R7�}�-���A �2\ע�"ч�mcb����(��c�,�� Y{ڇx��d	Jiʶ��,�H�r�
k����}&Z ���1�l��`L�,�o�^TA*H��'���������z_�����������^�E*�+AP����N��#T�(m��1������x6e�\b��<��x�rJ�B��(r%IQ�j*:k����*�f�4,30ٻ�э[�����>w�����#Jj�u�����������/̧����ݷ��7ꚟ��k���;س��?o8�o��9�A��$$�"Eɖ��xd{��Z�nMX�j�����c{e+X�H�"%&� �����p����ް����F޿�<U@u��o��9�y���~?߽�9q����\�|�cǎ��v�|�
o��6SSS�I��,X_[guu�����x�n�M���&�.YZ\e8���������q��nf�����1Nx��7�R033åSg�%Ug����:=�Z�|�,�	,�^x�,M�ENj�Y�!�26o�B]�x!8q�(��:~��`�*�Hcˊ���֢M�45B��B���s'�6��LԳB�u1�e`b#���h������5������RP�*x�����Kx�����q����Sϳ��h��;n`z�<hM��Ty��{���Pa����@ck��A�e�J�:��k���̩���Ͱi2��f�nߊ���8tCU��	"�Nc� ���qƓ�	�8�Bqeu�|}74�c2�c����ٹ�M�������o෴�z`J9d*�4@��6N"7/���\	V��rU�ٻ����\<w�×/�oj��4�"���!\c�
!+� ���OPЈ��KH��a�CGEU�hG]�$���<���l��sya��s3ت$�Z�a���o����*NK
[3.�q��f�n�DG�Z)EUS769k}@�^�M���QB���J������>�4�|��g�@��͛�p��/_f���,_��/���}{������3�1�ֆv���I�q2XЬk0���"JGAhZ�T�HGC�W�������d̖M��u�]<��\�r��.��~0hEG��K��曜9s��,��,���I�ƔA�50��*�:"��(�ÔÅ�=�?��-��"��gۮ]���甏h��Y�.^a���2�H��Ѩ?�?��PG�u��=UСq�h���跻q|Ō�������v���*��(��jq�m�s��Yևj�b�hl��Qĭ�:�-�I4��:�")IDg��=��Qi�|i�Z�t��r��)�g3|߃l߶!B��d8D���G?������~�+�K�n���`���:�ģ�|뭜9}�-��0�i3o��&gΜ��tB�E��4M�bM��"M]k�1�奫��o���B]�lݺ�{bR2.�e��6��5��x��cG9w�,�h�55q�C���Մf��1!j�6���fe�u�)�e�d<A��INY�l޵��v��'Op��Y�w�D�妭sL��9zf�������!�	���`�(!C�"� T�G��h�f/5��Aw��ԕ�b���
��毥]�®�(�fm�j#�@ ٹ�ۉ-���[��˔��������vmEZz�.Z*���2
��$\�c)$�Z0UDn!��z+��5�g�����S�5≁��kO�#R/ɢ@�[��6�u���(!��f��!.G��
eш�,EUP]\����c��/2�����x�3� �R�$YB�͐Ƃ�h���gc���1����$>x#����3�C���ګ<����K��g�s���4�EE$�ħ6��S�#@����$�S�$�Γ�+$�9��.{���ݍ5�<g}u���-<�v�ǖ�y����F���^���i|]A��<O�d��z��Af]��WIU�(�%I�AJMG���+D�>�>�sssx<ӳ���Ν>�357�z�O������i�����h�5!���5��A��i/�Lt!�t8˪�<��(����5��PR�n�w�4�fm}��x��{��㘲�x��a^z�%�^��x4
�k���{=�k�f���[�qoQr-�_����$��f!�BJjS��U�����D:���B Օ�X_Z�[[�W�}+k]u�]Q�E#��ϼ��\A�E�S�YgN�z��fo�2R����s3T�&"E:��R6�����,�`4f}8
`�8�*
��e-ULh7���8S���$ݔ�����ɫ1�RA;]3�X�ؑ70��O�SL�:k��m�^��`}���3��o�����_dǮ�����G_�����[o��ٳl۶��[�s��1.6�0�3�8�I҄����%%E^������2��$I(����[����ɺm���n���������c��S���g�������iM;I(�	{:^ya�D&���T�^��I��"�s"�����0g��Ct�g1uɑW_�֙���T�o��S�c��Z�&3��Z"[���cSR�"��P��Ґ��H!�#.-qrѝ��H!���TT>�ီD&��M�삑�h'P>x��8V&�Y�e���B� 4��;��x�O�<�?�ֻn�δ�lEj���;m�R�u�B]W�_!X�)��N�	������?Dl���Q�&:�8�ց��GA�"���-��Kle`*(�WKŎ�r���K��x��ϳq�<����)�~�?c����.L"�X&]l�HD���*b"���X1�}�~���܉Ў-�0k�K�����q�i�58j�v�����:_s6\�և��k�y��A�n�D$)y�`lݳ���̅�_D���3g��BG��߀��!iiZIX�yAKK�1({UUb�Gj�R��6�@���U]�G�\�)nپQ�~��3S���5z��m;���N �c~�&Ο�9{���(	S���)�S�?X;a{~p^HT��J��P��b4`8a��,KZYF�$��N��	�.��(e��}l۵�����Ν��w�cj��j�z�!�L���EKEQLȫ;�pc��7�M�t�"�f6S����0�K��u�w����p��U�4B�9n�
Fx�����i�6��2E������=W�A���[a���Nԩ�HVU���[���k�K��'1 ���S�}.^�H��b8	�pgU^��-����T�7Q�S33l��4�Y��^�KW�P"'�|���J���-��5���:��g������H!�N�p��96F�y�!��^�}�Y���w)ˊ�;���S����>���b2�޻�enf��G�kE�i3�K�h0f��*UUQ�V7�Q:��C7���M������i�b����n�Rc뒷_��/��d}�
_��戵Ɩ
�E��
��4w���k;���5tS'��D2��c�V�cV�c*/�����y��v��o����[�����U�.^D��&o������@��n�$��^�
�CU��N��^�,��Z=֌A��AYS�Y��W
��A<�h�5�9y��a�( R}Ho��Z1���૪+�O��~���^#֚��ϱ���q��qE:5�cf�Ϥ�W��~�o����f��S+Gjj09�b���c3���cޖh���6S��AQ�YT(h�4��ݢ;)���X��q58G�E��WT\8v�W��۸�u����C?�sL߸���I �0T)��Pq�B�P�4���JKք%޳��)��{���9}�4�>� �z�����o�Wӊ"�&q+�#�3D\K����߈V��?�Cz<�N�F�po�6$�u�fx���{�����
����L�zs ���o��ٳǉ�IYэclm�2�,�4�u�U+kQ�ޅ<wA������	�dL�5�W/A#���#o)�7�B�?E�S����`c��S'pU��-��V�=}��pL���I�X4�	�Z��>����1�Q� w��"�ʂ��H����N���fn~'���Cp�w1;�	c,'O���ǿ�h0d2S%��@x�\��T������%����*]S(E�5UYbk�D�J��GW�uiK֫!c[�Kǡ������|���8�w�{��e̅����F)��������HV
&E��*����s�9�U�$]OJcNYS�Q��^Z`��d�����H�	Ev�=��r�ݣ�iҰ����h�*$)k0V_Wtgi肽5�FC�R�qL�ت�9�d8@*E�fL����뇙��<���355Mv��U��K������������,�,�c�vN�:���
_��O1�i�SǏ�i�&y�7�����:a2�0u�g[*�715�%�"z�3�8fu}�N{����y�N��X��ȉw���s�pu�"�V��h�)���DM��o ��\'�5���6/K���t��Ye:aqu���;vr����K_�|H�o/~�n;��;�@]V��#\i!J�jO��y�8�:I-aU�wx�U�����c�qe��c�9VՈQ����N�<x7������8��+إ�t���g2)��D�@���Fx��)N�cv��Y�je����Ox��������Ͼ�;o�b���ٔ|�Ǚ߲#ć6�҇�����_)����N	&��̇�U܏���j��x+Aƈ�i���G��@�	�'������Hi����8 b����v�d"I7M���>�x���Iw�B;ƫo4$.$��*��]�#�����"F�6���RP��ʽ�}�����:�����O���?�~v�z'������+�
���r�qR��'h������犣aQ�0�Bb��F,Y�����-�8�ֻ`��F�?Jћ�q�]wr���Q��bIK��"�X�"M�%VB-���GX���f��隣F)��P�9��Q�ϻ����Ek�}����̢Zmn��6�ɘ�'�1.r�nEi���,-.�pq/�vpI�Fܪt �յi���-U]Q7D�k��J� �L�6mb��� ���ع�[o��[n���pȫ/��[o��������W.c�)�N����Ek�+8<R+�wTu�p<"��h28k���լSjo�x�2�#��yIḾC7��v����_%R���W^����U����N��L��w�T�U��8!�������+P����\A��%Q+��)uT��o����������w����.�l+��O�� i�ٵg/��i����tG@����h��FS��C`Rxjk���Q�t�G��,����E�겡7=M������,.^�(r��nv���7bme����?��o����4z�Q.^`uu���%�w����:��G���9~�8��ٻg/o����!a2)鵧p��?�%k'�o�D��E��v�`c8f����|��Dq¥�x�8��[��,3����+���(uY6� q	������uA�`m蘼sHcP�DE1VH�.�P˧{�5����y�W�ܧ>���E�<�&��ݍ(+\Q��,r�M�=�c�:��wf��A*
�JPJI!�=J[\^p)���������h��"TNv�^z7�/�ɕ+�UЖ߈��hv���R��)1
�:ִ�����t��_aEt�l#-{��ט߼��J���E�R�ˆ��A�4��`kJ�����2��E����m�� ��Ұ;55�Z�B+��X�b�C�����A`�]�U�Vh��E�~��I�-��!j��b��s���pN!�-H=>L0l��̙��������[]ض���ѹ�v֭a|�����O<�K_�S��5n�����^.|㻬�U(�Y�j�N	Ls�q?ܡ#��L#�3"xн��&o���I�eI��L;�N��L��B�"�����'Jc��~��RLTF2�sR�
��kЖĻP�Q������&�ܽ�Ml�$�B���o-�%B	�/����c�1�{�gמݴ�mn��V�+9q<��&�$c����S��}��W�H7/���P�l���m8�q�@�ŵZ-�4%�#6�o"IS�6h�����[o�ҥKԕeaa���|���:Y�r��e�|��j6��273��"������h�"r��E
�3C���GU;
[`� 1��T^�H�������I�������s|�c�VY>z���U��[Of:�Fp����(ƷہI���s�������_��(�֑��9��ʆ�o�����ѣ��f�M�TUAiZA�;����[n��_Ak�������T����2���~/�"p�M]QWU���v���I���1de0d�[��t���˜W^�>�_}��}�c:t���)�k-l�XY_��e�ܵ�$�Y_[���ؾ���,��v��烈0uM�ףߛ���e��dfv�v7�b������ty�����w��-ۨ-����>s�4MX[[���3�k=�i�O����Q�I��N�1bmr�,�Ѝ^.�.�P�cj���Y�IU �����}�8q�8��;����[��y��B�1A鄢���0E��ہ[_��������BҖ�G�C�7R�ѻ��H��1I�u/��ݿI��A��)_8�ڬb����}�'�-������::Q(�F\D��uR`J��y9��B��y���M����w��c�ƀn��K�&��R���o"���%�S�j�D*Ǵ��#���?b��w�5�cJKRoI�.�P\q��� {ￓm;wr2˨�
�c<�TM�@`�ǣ��N4Jk��^ff8�֎�fRn����TY�T�}ʚqtM�JT��L&D�DF].l�Iϭ��;�c����ɸ��>�9��N��'x�W�����;u�5g�n����eړ�$m�6��P����1�טqM�rӭ7,wD�x�%��L�'�h�k\>v�[��(6V����ܽ�{��g�z��9j&O�5�J"��:4 {"�5���Ӷ&pכ�kj6��A�f�U�SӴ[]l1�7_c0��{�e����=�����`��Ǐ�1���%�2��?���-,//�1RKU!YQVDy^��,V�4Mhw��ZY`���t��6o���}��t��&N;��j��n�q�q������T�N�������qW*��<!�DJfgg��6T�^��k&�A��H��ݲ�|Xr���ؾs/���<����Me�������F����L�Y�g���&��IBG�!}{��s©�\�jh�����ʺ�on0W�Dy�]ҝ[hm�fX���A���;����ޤX*���(�{��1&ؚ�$��f���4U$Z0v��T[�T�B(M+R$qLe-������������y���_f���lݶ���5fffH��K�.1�L���4afn��-�i�Z�{=�9ʛo����>�7�ȱ�GY]]e���z�mL�O��p��Kɫ�-33s�ۿ�V��ٳ8|���b����gO�`4�`��A�%Y�`�c,��P�B�콠��������!��Z�)$ց0e-2K�
O�n���M�?�g�x���U>���S��\8y���}��s��gY]��r���Hq�RVJ"T؝��E]je����H���2&���4��_����7W����댏^d��8�����_�"7~���Q���CzA�@7t@%$��R"<3:E�T�+-����Wjb���i�ra�zuHo�ؐ+���y�����oﱉF�"��S�����u�2���KW971�����qL{f�V���J��,��(��PV��$�1��1B���,��R��x�?���p��ɹI��.�ׂ%c���#|�÷����	_V��"���
�8E"y�g�硻�ݲ�=�!���wy������
�.��g_��k>����=��'�ͻ�M�m �9W��݀e�5�א�PM��7��3��y��څ��#�� �������K*��4��&k��}��~�eFk+�2,��z*a�6�k�78��ì��8��Q1|�`e��R!�Z�qT�!Y335ä6}��=~��{�p߃�s��*[s���Q����cTX���i���ͅ8�IQ`���ig��&B"��*S1O����J����o&JSV�ֹru�|0����|<fzz�b2��sZ�s3��UM^�GC��"�1Z�Dq�x<	�%�t�2�V;LO�{^4�:��<��D����D�C7�Nwz�^x�c'���?�c����%���Zb��ۭ�y��aEU)|cT��}/]�ɂn��*�I4����갎�;eU훳:�x�8�-���¥�Uf���c-���϶��9s�4Y�!��
��E�2=��&I��ˊv�ZY�R��5xkɲ�{*�I�������X^��S���n����p�<�������(�y�&�	��e>���diFY�L�v��h��淾͖�yz�)���N��ʕ%��D�f0�@G��� �e]����	��o��2Z����R�,]Y��Gt[)�;��-�Y�����A^V������P���濅�66,�B�����o��ɓ'�r�nn��^}�q��9��[\=y��pȦ�EWǴ��:�� 9<��*��=�;�4��S0B�I�&���"F�����1=��]�o�؛��W�1G�����qS۶����I3�bBj�[���c��	��1�
V�L����G��:�V���D��.��A5�����?LXQSi������>�Z	�3�T�t��>���A������X<~������G?Lr��%�e`�K�<�&�[J!�(r���DSG
3����4a��m|����*-i�]s�O�������|����N�K��d��D#�DG	�:?������s�w��|����o���*�d�L&L:��?��>p+~&fg>���o�qd)g�[�B��&�c��&��f�n�p#�Ct@� �HS8�h4b��9N��6{{)r�*S�=D�f��}�ڽ���W�R�ka2�y�	{`�$�$����J��k��:t�B��D)�����z����4���xȻG�pu�*�n����(Ŧ�[(�C��#�1Ƅ�FߤJ!QZ���?(�B`+�x�SU5���[��{ `��m����*��o�C��enf�a]��(�Y^_��i���N+Kپ}[X�yO��c8 �'�b�	x�(
�1�5��qMڥsX�K��$Q�H}��	+W��s�F�tgϜ��_c�έܳ����\9�.:�!i����R��^\���u��'��ɿ��_��^�ɂ�w���'���{�,F����X�8���p��8�ڼ�pQ�����l�Nq��%v�؎V�4kq�}��K/7�r�1U�;��aye��,P�琑���FG�8���12$iB�Ds��x/X^[Gǆ����T��h%Rq4$�Rʲd���u��p���+l޴	�,gϝcfz�V�5�Ȳ��^"֐�%��i�����3H�kv��I�,^]����Dq�$m��2ƃ��P�c�3�{�صLM]UD*�"��B��آ
�A��Z�¸ ��>�3���X]Z�;�g���;mΟ?GYL��� __�ҩ���)��g6$eI/���I�KR)H�
;�8�n�Q�hR� -��d"e�HZ[w!�l��`����;<��D�6�����m.=���zI���3E�C[;���"���v��T�0.�������E��L�t�B��X3�x�\$(�������_�W#2Rx�.]U0��I�g��:s�s������̿�v}�S��ۨښ(/)�#��t�Q�(�	D��)��7�"��*�n��d}�����[�.pŘ�_�*G��7o��c�G?�q����T�*iӲ�,6h�|yg��{���8��������{�oA^ӿq>�[?r/�$�#��t�����z:I��QUg�a�B�j!BA�a}��20�RQ[y"U���L]��x���%V�%��#nelߺ�C���[�3�������
[�h��2%����� j����u!��`�o\`���ˋ�eE���ﴹ���¹kkk8�9t�M��o���~!)�k=u�kki�ژ�!�F�?)gƘp���Q�&/� f��$���a4�i�Α�TTL&�9y�V+e���!X�r��Q�I�k����<P��{GU��q:v�SZijS3.r��,FiV�WȒ.w�� SSS����//��O���9w�]����ad]�;�kƋ���
E�V�͒k�����,�����kl%'���,K?�Q��bP�G�Һ���ge��hأ�N�:�ƛo�я|����8Z��/�Y�2xW�֩S�.�䢘N�G�O��DQ�NR�I���^[��1�$�=&�Y)��9�hcH��F���*�Cʪbuu5$�W��n����'!�@ B~�E������Ī5�,Y\\bvv.d6��Ms���1X[	�5Q�iHuJ/M��P�ec
"�E��B����"R8�1XSSՆ��x)Q��<T�"IR`�g۶m�NO��K/1��r�7�ړOa�7h�5qe�Ƃ�T�Ȉ)�h�iy���R7��Aa/]HM�|@�:�Pi�%eelHw�f�C>pѹs<��'y�O��g#�4��?�[�S��}+��Zƒ"�?����N���$�ᑞޮܿ��7Fj����2l� r�8(�U}���FJ�^�i���|��J�T�F\������?e�|�{}����D�民FE
a�4$�%8D����o�>B���AF�,�q&��Q���.k�p�����է�`��}��c�b궛�Yk�J��؇`"T(�Z
TY�s�<�(_f8^撯��ٟA��̖$[f���>����nk�hLRE�~�]�Gn�
�~}��dBK%$�"���C��X�܊ƛ�DIE�jjo�N�9DU�|DGk�u��5�$f��D�;����:p�V+���՗^���s���#�F	�u׆Y�������
�cJ��j������	:�C'���yQ��;�O�k�k����(H��CH���v���!EQ�n���:�h4��*��4�1�QOj@`�a8�"(Ϝf�֭��m�<����s�f\m�:Y!�^���U�"�4E�X__gvnk-�ᄺ6����ֆC�T����N�����pHa�bL�<q�lE#�  �5IDATa�����}~�u�x���ζ9�i�b�
o�җQt9��o��]�:�.����I����]�޳}��[>��y�֧:i�����;������z�M;�1������n!�t{�yם���k�ҘHJƣ!uY�RO�$�XhB;�ҝ�AA>P�:�� �0��&9B,d��EIEY��b<ɩ�1���׌	A/JSYC'�iE�D��bem-d	k�����4|Hw�.x8���H17;��>d��Zx㘛�a�?�x4fy�*xOQU�c�l+%M�s�U��\�G;k1j�um)��HB�P8�]MQv��Ida��Fj^^�q���Y��s��O��S��w_{�n]�6��L{I��9G�C[�N�L,b|c�އ��������4C��b���]ZY�]<�c�O��Wac�ݟ�$�M}v��[MX�ַ��[m������)��CdAD1k�f$k��;�ܥh��j�kCE8D�["����ݘ���/"�DY:#놕?�s.>�,�%�Oui�	�ç)^;ƒ���~[6on��:�8&�}F��D��B�S���fb5=#���ْ��_�ԟ?����Ю����O�w�EX���r�t��AAjwx[�|M7��l�xX����\����S݈�~�S����+x���8�}[���#��;���'im���ɧ���ST֐K_�Dރ	E�&�OyBJh��R"�_inQ�&�0�ns��UZ�ӑ����.\fzz���,���ngy�2���☪�I[)�&���F��okey��v���Z�y���\Z�����`R�d�0����uY�YY+�j�Q�ᬮuUa��(J��)�I�R�u�T�Q��@���hɌ��:�l"�ӔN�CY�7֙L&Dƃ!���5�,���zE�p8hn\���v'c4R�e`T�մ	���ڗqp����;�����bfj��K�<�ҳ\�z�?�)�ӄ�����cghՒ�ɸ��>�L��SN��G.I k�j����-W����{��������/����J3l4�V��4�qߎj���L�D,���o�}��^��pХ���1{����o��g�K��"��+�aUưs0��F�pUA�":�>u^ଥ����qJ�n�E	Ic*��`@5�1�"�DZ�	����pB��1�vF�ݢ,+:�6W._i��	q;���`3�)5>� �+y��cd�`	ٴi;��@I��=y�Օe���LϠ��Et�o�d���MGQ8,\�xj�1LL(��f|C뺆��\ǡ;���"�\��ٵ6Mu��G���)V���Z��gJ(Z��i�Z��I�$2��T�zMP�|�m7�h�J3�Ă�֛زc/o~�s_�w	͎�`��;y`e�'���0��ܧInރ�s�gX��7魭�f�:Åk�/��2x�#�ؖ�H�[m��w^���E��6��M�X�E��b��A$(	���0��9;^�`�6@Ljdi��,���!��ޭ��W^z��k/Q����)�w��25�!=(B��	B��%�I�	eZHD���6`���җ��:�i#aa���<�?}�f��Y�=���S�z��NrMTm�ER2%$�ڐ��Øn��?H{�NX[��ˠ��t�CC��}{�� #@ܿ}p��
Kq��fZ
�*�:ҡ	D@�r�G ~�^�ki=X��=֊��x��yA��p��w�s�6�$gfz��_~����ȶ=��ȇ�̱�\��n���)��X�R�0_��a�_�=�P�X��]7���yTgF]#�@kA�o���p}�fU����l���2;է����r�"/�w{Tu��g��ź����v7fvnc-�^�~�O��1���n�@�R#���XQ�$	�yb�)��Ԇ�`@U�(�H�ck��0��M�Ir�!�b����=���6����P ^򢦓tعy;{w��[��6GO��m����Mq�W^{6JF��u�\p�/W5W\���"|������ם�{��T��B�Q��F��Z�7�VWn��[�s�v������4�h<"�R�$��v�m���˔�	Y�P�[MZN�Bi�E���v�����&/�O(MI��+���v���B	�`4&�*
c�i�hR��"R
[[�4KH[)UY��O155���4+K˴[6�m����x�tDYV�8&R��>33s�iL9�9{�4�$f���.�ne��{�#A�աGS3O�&��Q������	�'�J�ЭM���=HH��9JG�G�A4�H�8�Q����O~�'8w�o���8"���:�Rch�XE�h���l^�^���˦�7�w+E�1��l��#tn���o��g�������Hi����롻x�p���~��~��9���3:��_���	[��j�L�����Ip/0e�Lb"�`�c�V�8Λ/>��7����y�Cd;v���B�(��	��N%�RT�iIA� %��}<�!*r��(�Fm�Li��ۑq�P
-$�"2�ktPe����C�� F)���ҋAjA���t�tt[O8w���"sw����=�qN&!�+�C"��҄�'����n3���"����r�Ͼ�}��q�(Bm����?H�l�9����ʋl?��-[7��8��Kؤ$�D�+�jg4
�%��OJ��8��$��8/i��3o���&�K��m-�^����j�8t���~��p���I�S�$:��BzYar���g��agEmT�w�D8�]�pֆ��TD�$�ઊ8���7P��k�PR�(�T������`4�è]�,�̄t���A�n*&��4KP�g��(�P�-�n�����p��p\Xo��)i����(��4K�qD51!0��@;����s偼ȩ���2l�α�n.�9Ûﾁl��ﻏn�8������*�F�'����*��*e���,�w�X�~v��/�������+��/�;���*#��n%����3)k���1�M�3���z�*�ػ+��n��V��N�~�;�J�5Z�0�u��W�"pL��XyQⅤߟ@H��I�y���w{�Z�@b�ֆCO(ʊ,I�EI]U���qޱ�����Z������n�صkE^��[lٲ���H��v���˗#�m�J]�,--S�'�e��S�M��u;t��n��i�"�k�l��^�C^�L������Q�klC�	�@3�x�~�k/�~��N;���=p?_��_e��ΦV�����'C2��t�D+"ʂ��z�s2��h�>��o+�2��
;�t��1���ܛ�x����O>K�M�y�mz�!2Q�淾�����s��6����m��V��Y�E\�p��>(��݄Qe�Z��yx�#��:ϙ��[O=��7/�����}ۭD;��|ш��Y֚�/���������W@?e�G��`+�j��^���
�#�
��&�B�h��D�wΰ�J��sL�Yg'w��_��x	Q�A{�
�}rю혖D�N��.� 'C(��n���Gb�8#t�R-��.~���6��L�]��J�q,|����3��n�֟�	ff�>������R��b�uR��sh�0�X����5q�)'���v:��9�GD��mܰ� /��&/>�<�=�0�<�(���»���B�(�*�H�]�c�&�A�k��*�F��7Ht)�h�4H�4���V���25=Ö�۸�x��h�0IJ��ƭ;��ٌ��"/q�S����|2BȐ�0h��3S�#�#R�|�+I+k����REQ�|��)��{��7��!�0��Ĕ)�n�4\P2D�BP��G䮦?�g﮽�u�y���Q�྇����t��'NQ_]A�Nw[ozėk�Wl��#��w���q���,3�Q]��0�T��[)�.\���4m}ye#�=�%���
g�~�M7d�����k�]�����Moz�䣜={�3�Ob�Cy,Y��Z�RA|V&	Y���*W��v�g<.�	
���E��g)�&���0.K�k�ZS��$&�!ڢ`c�#�`��a�ř���{Z�6/_��C�H����
~n�ŋ Q�V�Ic��5��L��`-�d��e�,QxTa��r)��IY2.+��QYO�<������D�Jv����Z�!VZyTS�5f�s�7�s_�<'�x�S�_c6�h9K[B&��L��t����U��aʁn^�J�W'DqbL�B��[()>�F	������<6��'��o����M�j��ݸ���Ǖ�G=ɎR0��)q�aT&�u���
�'��D(l�C,m����L��̮��b��78��i�<���*���^��1�"D���,�P�>pփ�yJ��%�v�d14%Y�B��`Y�rԤD�u�Q�v��*�(��j�^~�w�ދ�%�b�Hc�3�o�Ǫ�H����;I�@ʚ�T- ��c=FI�އ0�F��6���FJj�)��e
�<>�U?X��k�;-���D��U��^����v�>���0up���>�i�M�9�����י�"�38߄�8�4��!I)�pDB�Фi_Ԭm�O��±<S--q��	ny߃L�3����s��"?��?��?��t�t���H��>��'��f��j�ıփl�
��1��a4d�bD���g���i�@)��f��4�~SUkI#�s�r2&�4�l,� �n��z;���G#���鴻��8�`��n�ME$J3���v�ֈ�V��h4�9G�DXR[Y���XY]F)lqyM��Q:�^lcˬ�EyE�8k�c*�9�VƶM�ɢ�'O��l۾��ﾋh2������<�ݘ��R�n}yd�׽R�F�J��a�{�v��#P��/���Ư�� �.&�<CkݷlG���?�Ս���\�����3?ǁ�;x��1�js��8p�<�������?cTl��ZĀ-K\]�tbʲ�C]�tzLkk+LOO�u���^P��xL<!��QU����q�(���:l�S��d}c����)QJ�����%m�XYY!�c�[6s��ƣ��~
[��̄��Ob�%�*.=Ji��S�nP�����!��-�)1��ـ�t��x�RQ+(m͸((JCQՔ�am�O�BR#�O�Dy��iEaY�0��n�LA�ӭ6��s?ǜ���}�ykٜĴ뚶�d
���ј���q��I��"�5�YdU�'9�����)�JbZ�Ť�,X�.��(���[���s<������or����.r�]^�#��M�� �I��fC�׺�0��z2W��%l{#��dF�����y�=�ʱ?�3N���]>������;�B#U��F�qtR:�4!6B��!�E�A��	u�CY���S:Y�����2���������s��~�t�V���T�ҕ�6�x��X~�ʩ�HW%� '�y��r�2���l�a?��QJ���E���6Õ!�����j�ؒ�DHL]Bⱦ&�&L9�@��yOZM��J�T>gZI��
��qʹ^����S�n���?���vr�ݣ����L��}p��|W԰���:��Β��9���ţ� _�emT�LLA�Dt�d��	�7�0�:˭�w��t�ǟ��~��x�[；#���t�EQ9t֡,FX��l�AK ���;;��$��	{�8��q�u�ڕ�e�%i�3YP������,QZ#����!A�*I����#�L�X]E�%sIJR�X3h͎�^�5&xO1�SN
ʲ�x��./p�ҡP�I��h�ho2 8d�V�t��,(��k�P� ӝ�$)����	^J�Ɍ;z3���9~�<����{?�}�r��?��S��q:��g{O�|�P�����)�R������C����|A�j��S�Vg��w4A|i�,�]}�Ta���o�v��և���x���ĝ6[�m����ϻ�N������dLU���8�KO��M��G��&.˒DG�J�[�4�s!X][��jjc���5B�H��m2��)���.x�'EIK*L�� �i��ޑ���UI�#����T
6�o&�
���Ɉ�b2�]��2$i�:�ֽ��u8�KI��������:��;�/J8@B���,��Ͱ12���� ��'�D����о=|���S��ϳEk:eI_G(,��H0Z�j���8N0�g�r��H�"�#R�`K�n���%��]tn8ȸ��ϖn�h���v�\p����|��C{���|�7��y�~�}3S�ʜ��w�&�a�}�����h�FV!�$G&m��a�G�^����E�/��d�ܶ�d�4���.���2�	�6��E�hDx Nidq	�h�F���_af�N��~��2�ΰ{�>�N�f��#T�|�t��ٜ<�
�?'އ������C��X�ĕ�����ϼ@�[�a��c��gim���#�񹅪����F��D��5S��`��#�hho �%mS15,��̦V*ËO<C{�Ã_�"���L���W�������l�e/�w��駾K<�Y�x���DD$e&�X��k�TD^"�d2a�����@hA,4�1,=�����2�>� '/���'g������ÇY����EU��Bs����?OJ4�JR[�c�k"N�Մ֮���eHoA.a��(���5�kbZ��`L��zO�AX�����>&�1!D�����˚2/�m��cjCm-Z% ��+�&�cl�>O&�Ű�����Ҡ�a����M�q;��Ҍb��Q�1DIL�"�\]du8���e~�_�w�ť^��w_įL�2�������+uU��"rBG�v�n���{���(����?�k���{}���/�w��g��k�+;6Oo��Fc����m��`+�_�֟rϝ�r�����G?����s�mZ��=EY5��eQ��g��qPr�/u oiB�0�*&�1��$�L���T�Bx���,I�_YHjg)�%MZi�VZ2��PUZI:�6�.U���e(���7���"�2пL�P��N#��"Pބ�xCU;��`����z��yӌbL�H*hT�!�9/ ��%E]��ZT�P�!R��[o��쓼��'8��6�:t����B�ֈ�*o�h�������A�K����:&w�{��1��;��g�H�����NA�@��a<���O �=�]w�K�j�{���w�bM�5��� �������î2��ә ��R�R=��s��#�y�5.?����m�ֿ�f�	�e �T���7*��5[\�Rta����%K����?���F{f���`�'�����}�c�?�����=(��0]����o
��+U1�vP:dQeH뚩4!?�o�����'>���3�ח�X&��5�M�nP�k��F4 	�H��)�A�(��33�,>�Ջ,h��[o���=F�L^;Ι���W��-+VN�g�M{�4�	�%�&�2�7 �wO�E�vlU!-D��w`E�'0��;f����r������&����>���֗��'���y7��v'�a��e��um@��/.�O�yN|HbS*L\�(f!%� �TR4x۠R"�\s0��j�U���s���û@���Ǵ���Tu�d<&�!�5Ѷ!�4�pMN�!.���P��`�$E��/y�wa��
U�)d�	"E�$DD]�Ԕ�;���9	�4R�	�*�,M68p�n>�鏣Y���O\�Y����t盹���Pz��n������?���s�)� Um�q��v��z���]�Iֹ�jQ?2Eڜ=��sϰ{ۏq�]���k|������
�|�Q~�S�q���eNwz���:�8�[I�WDR	I�+R� �;=8`/��dI6�z�����XKI�΄U�����)��%�Z6���<��^!�ݘ[b���0%��p@>#D�:�^P�%(�$�9j�Kj�1X'C���X���9���k�uyH7+��(I@*�b}}�=;��~�?a�p�o�ᗘ�/�Y����xO��LgKÒ�,0J���J)J�P�IA=;ź��_]��v��4�0����L�kv���x�I.��-!Ξb�Wt������p.����Z5��*�����bd�`�_�����_�3�$������>���;��z0�b�A{��+L!����f�.�'ÈzdH���a�	�(9�7�t3Y#�)i�!�g�=��+�}(4�����ڦ˪\pn�����ի�+�눔f��I�C��"�+�P�P
Fe�`2�%C♗����ʵ6]xP�s�<XZSՠ\S��u-�0��������J��8u�MN�?B7�`2AwSbť0e���<Ǌ�R@eFkV���m��I�TDH��#�l:Y��R����x��'�S�k��������������G�5���;3�x8`c2��~y]a�kk-Bb���5a<>��e��k�G�w�(��u
�B���*4�!T#��6���HEc�X���] ݄��`?+�������p��3%��(C�ցt9��!�^+<M�Le0�
��H�p��=D*j�piCP�rat�'N4I�����L?��_`W;��w��>~�VRU�f�^����ښ�NkO�঺�iD�c����������'~��_Q���1ea*#g��o^��t0���jȕ_��c��G�O}��ϯ�&_����U��?�A>�я�o�)�����$�C Im�J�xF!�N�{�k\�@+E���N����� �����k��b1.�آ$�4c��QC�����D8��aklY�j�s5I���$�,��N�q��0_�;���u�	)R6�����e��a|�ҝ́ Pٔ�+�=� 
r��	VHƓ1���V��7��/0�=���~��1�[�kcf�U��F$�Z)u�hr�b@�3�֛���X�cD�4��5��U�7r�����?�Ο�f���S�E+����?�]z��[�`��e��++�|B�-��C�4
��k7�����V=����٦���fU]�˂���8���}�S��M{�4����[Vh��))��v�DJDx�f����.�]�ʰQMh��V[15?ťw�fϳ/0�Aа��1�y�0�N�׀���nʃ��kbFD`�#���Ւ����L�^et�2÷�&�Xb�*Y}�U.�w�3Q�To*�*�0%F�$�� �>)Iʆ�\*I�<N� �]�jK��"�_�-/"lf�����C,����w���G�.��x�5�ш�$f�����X-I�������ZC1�mY\\�Si�HxZZ��,-��@�tĪ1\9�S�q�g���8��}���Ffff�z]N�8���s�2웅(�@x�h%�Z�p(�|,��E�
�»#$@
����=���9���("����n����|m�x^���TS����p��lS��D �B����3:rM%L�ʔ �EIm:���i�R�{PR�&$�	U]!�'i�S[JYRKCQֈf�eK���*�?�����������c�ר/\����H��ۿ6�ʷ�R��Q���X	����{��?��G���&9�VJ��`�9��t���33�擟Ͱ]6V9�ēt6m���w��?�~�7��}��DI�m7���x���9̠����1כ�.'T��5
I"ƃsdq���Z�)����'�#���e�p��u�p
�l�V�s�qu����AJI�|�<B�H����F�	��8�(!��НY�*�(*C^CY[�2A�c|��;9F�H�9��6|OB*T�ZԦ��0U�O�[|�'?�]�������ƙ�iw���hM\TPVX���Ś��)2͖�o�·fz�v���[lP�!A��X����S��Ԟ3�.���|l\s�g>G{�&�2��W^f[Y��CO����I��Y[�]�k�:\����\����Y/
.鄃*gz������q?�����*I�f�g�$QU��+��Q��%]���O6グPB!]MnGTf��lĭ�������������|ͥ+�֗y������������c~v��I/�͗�!S��,�uŞvB������7��$Jy�k�/r��gI
8x�}k��
���hH�N�X"�������@4��dEHpvaHi"N�Y�y�)t�Į�������܁�J�
I��8���8���dUM4?E���vK�m�j��P��,t��1�ᘅ��x����0H�0�Wޣ�#�2��X�X9q�A9Fe1x�Vk~�[�d����F�N��D:Vk�����j�F�(��AU�$IP�Zۧ)r�yDt-��7�� �c<��(/I]WEI'��`F:��L��A]4L���=~mj�k!�"����9��4^"��l��$��2L�T�$ت��PI��γ1�PYKm�N�$k��D*�g~���g�8���<���O&���{_���I���V�i���Ri�������G�������W���%2k����!%�i�JQO����X_%����ڷ�_Kn��V~������W�Ο�;o��[��r>`m�����RiE9Z��je]��`��*���[������1It��:K�ݢ*K&�$�^lB
�!2�������x�Y�j�݆`g�֣��T�!^Tk���6O�n��qi)j�{mA\pИ�P[���9h�f���N�v�����)&L�18G��}��|�������W\8�*;��NQ�
"+𹥝eL��f	�Dp��?���=�P�ӫK�N��n��aT�e1��twm���)\n�߱�7�<�����8��?�I>��g8�J�x�q�<G�I(lux�*��L}m,��_ޅ�B� �Y��X)|5FW�+�G9g.��S�CLr���;��t�mw�Bo�۶�c�#�xL�½SE�����?�6�w��c2a�k��e*]�̱V��/0�377˾����N0�s;��DHQ��D�0bn���y�{��,�p#�Z���,&�uniŒTxfz)��-Y\����9�he�5y	-��B#��>��z�C�dx�1�QaID�0��Hq�#\�����O��Ī����_�:��y���
;��d��w�Yi;&-��QU;G��LD���9v�N���r��ì/,�6�'��������m����UF�[->��Y��Ή��$���RNrT]��)��X��(�ъ�E�p�ёϱu�-kUU6�V��R^�K����&��|٬GB�G��a�����i�4EiMU�k���3w�z�~�ٮ����`5mv��A���I���ֆ����^ =@]��d��G���,B���)�EE�N�ȇ?�O}�3���9��s��{�!Ϣ	Y�D-��8ǚ�Ÿ^�na��y�����#U���?����?�ȩ)�Q���*k��ڭ_�*;�<ݿ)�N6���l�y�m���[�6� O}��y���d�M7s�=��%g����*q$�[i���`�eI�$q2���FI��*�	�F�T�nrS�d�5���	2	)/�"4�5��e�᤭d8�ΣP��[eUQۊ�t?$|j^�Γ��IY��������o��6��DO������!k�Z3�'#6�W�����?��~��9��wy����!��$�J�����hg)���ZQD�j���G��'��,-RH��$�Wx�%5�Q�A�&�zՊx����������>v8D��Ө"'���%��ԃ&� ��1���e{M��EH���	�n�������o�αwY�ؠ����`�,�P|�;t�m��^�c�q�������*��e��x!Zध�0ɇ�Ƽ��a_y����iϝ�����,3�u�L��7�ϴ���l*+��(��+ʪ"u!qL�0j^`��ҘpBt{�"o]����_��5"���025>��4&�{,�Vy����(W�tƓ�4M(��f��D���^ #MǮh>{��"�ㅨ頙/����D[7��]�N]��K������}�lG�sn�E1����Udh
%1J�1X�Z]#%twme��w�k,_\D�(�X�ڔ�QBTUd³r�"[��v�Kk��O>�)ʯ�)Ͽ�=c�����u��[�4y�IA�d�ZQV��q�"���HIe,�ɛ�8�_m��VT5./$s��Y����S?"Qui�#�L!B�tUWA��(�]��b7G�Mw�t�=��˦I�G��p E���. �D	�Px-&�����EjAm4�>�~��O���O>��;'��e佉���U�jQ��Nh�ƦLMQ��O����r���#W�~����?�/�S��U���)��eIkn�^a�51B]~�(����>��M2�����2���"��&��̉�Q���Yd�QN%a�$<�p$Nh�����(������y��t#�`	�p���ZE�d�j�=k�1�'X�+c�mȆv�����yYSV%Um)�FP�𒭽��*�
��ׄ1B4�[��-:��OM3���u�-
:Zq��7��������y��])�"�Ɍ�%t�X����q��������Or��k+D�&�a�o=�Y, ���Bz"Q�s���A�╯���n���U����Sb�5��k*�5�TSQ��%x�s!4ֹ���؞�"���7F	��l�5Gw~�,��nwѝ6�ʰzy���Wy����&%���Xꢦ6�Zt3�p����A9F(�ܘp�W��?Gw~��&�o��{�وD&tJ�^:��KW8�g��Oj�e�l������چ�'�kK^x$S�.c[q�;����X��E��0�ψ�L�TIL�ju�ɓǱWW��ߣ�i��[C��6%^�L�C��uH�C4��i<�U�_YG�A&����c��K��طs+'�;?�:��qer�������*�$X�6������"D�
`z�6n֊��y���!�N�rR�:��;Z�/J��D,��c�vV.q�������I^���7h��I�7�xc�d�ϴt��<U֣c�NZa�U�
{!���2��e��� 5�8���8��\`���	��T�H�r����Ĺ.t�Ƅ��\3j�xc=�7M$R
L#l��Q�f$a�sa���oq!%xk�B��?�)�Q;a}}��}/?�S?��Vʱo}�w�y�Τ�2��Qz.J��˫��Y�Hb�?գR�_�_~��9��t�g��b�Z/�Y/+���&5�(�~?����3/�H)J�������B��G_������LMM��3�VF�l��im&�uP�`�S�q�����$m5��A��5�N?����u"��`km8$8}�l!������恳�c���Y��Z"����,�Kd�Q�����8!�� J)���Ԯ|Hwl��TuEk�,���C�����#�Ϝ��~��L疸�LH���b�%��Q{ﾋ��Y�X�����>�xB�m��(���Z��=��A�<k�����[�!/�r���<�f����F�)	BT�b.��o���vF��	��ꚢ����ɤ_�'�<ȝwޅ�5�F?f��`j��QIB���M�ܢnb}e���N�q�$�T2�-2h�6��)pJ��ab
�&c�N�����}�Ѧ)�vn��R�.�L���GCH3n����q4a����:���q��p�-:t��2.+jQ�P#0uͥ�'���;�ڳ���ПjQW#�𴒈�ڃͭ>��5,x�ǹx�2{�=�Qܡ0E�U��8wP� ��<DΣ<��B�|]W�{O$�NPiL]W��i*s�����u��\X:�j1�J&7�:�g��PyGeU��֣�h<т�Y��)n��C{�yVr�l'BK'��W&t�^��^d�O�N�ks����p#��o������q�������X��q^k�V�V�1.JFŀ^�Kܞ�W%��Cx�c�P؃�M���5>P���$%NR�y�iDnR
�HQՁ}F�ͺ�r��\�kq��i�mW�ـ��JǁF�]`ox\�����Y�U��m��!J+<�)��D�C�������ʮ~�7��Uο�rR�>,�����o��#S}�
֝V�,��f��я�������G��������!�XA����N���c�~qei��n�u�Gډ�j�-�~��y7���_{����cg�1�%ISu>bS����M$��`i�;I��D�G
���<���h7�!\���sM�2���M6�k"T��t]U5EY�]�o���KU���"P:b\TL򜢮��m^�_8D�	�BJ�R���y�>tL�O����� �o�u��r��gٙ�N�e���dkC��Bk�~�e[������~��,C�-]!�w.�,C�Icwr��k�H4�Z�b�S�97�8����+��5fK�.��/]�$
$��'������҇ĉ��R��`c4
^y�0N��������G�8Xa!�\vc�D��cڥ�DF��u�N��me�ф��e�W���&5iY�U�N��eU��d�(�u�����L�{;�] ������,R��z��SxI25�ʇ̘
����;G=����X^gSܢ�S�(�*-�#j+�����恿�y��.k�PǎH9��`�ԚA]�fQ�������۸��˼�0�/��&�s�ҏZJ ]��%B{*����N��C�qRs��[�`��e�����
$-K˹,�'�ۿ�zKq��;ĉ���0 i%('%�v����xb�6x�KW#TH6�8�\p�[O�V�lQS���Q�T���4������}j�N.�%�|�c�M
~�~��ϱy�V�T�1k++�y���MH)p�1���I�����`A�a�G	:��Mf@YVXc���i����·�y�#��e3Z�V�!�A��vk]x�t2&R�0j���3K����{"r~ ��F�/E��ckb��P��aP��RkGU|��>�vt��������\�J֙�+K۷o��n�[�R8�%��)��)*)�����忕��o׏l�0�s:Y���p�ek���p��Nsz}q�o�M�N�H,>������Os�#�����wy���c"@x���u1a��oBD4BEH�p�3X�iO�&h�Cao�FU��i6t-�5�	;0�C��u��8D0���#��x)02t�R)�2�V=�0)k�"D"�1�ŧ�&���0�nF�צ��.�(��vyy�ٙ)���|��|�Ü�U^{�����e|���6r��f\�x�(�c�.�~�����gy����gHfz,ש���`,�TdQB+���Ck�k��=�����U�����c6&�Rɘ�4��2h'�u+�������>����05���$9��5�}����/p��i6FC�T�� jK13��j!������Ѷd�}�١�I7�;G�&ш$@ I��I�� ͒%Q�����%-{ylӶG�cqdk,�$��(yLR�� �HD�FGt������|b���o��uν4��@�$������[��N��/}Խ��tB_)�x����>���MdI�\5��::���Ԛ3|�� �ܺB���C�����Q�2��'y�D ��A�Z:Ǘy������֋�X�$Ld�ƚ&okWsc����%�q�W.�@zd�����=���8OUTt+t{}��cʺ������џ�#|��W��<�NPN�w�������Ķ�(�zp����NYT�\�!��%0�3�����'y�����"���M���r�N,X�t4fog�X��S���ʀF���w����җ��lZ�f,)��IY#!	�ᰤ�$�<�~wȳ����%��g~���S����Oy�'X]^����̦3ʢf{8$K3z���3�gq���j*C�egI�L04���yp�xn>
v.��2x/��3)fM�M�����_k��b�6�'�n�a�m�nM�UT����}��>
 J�"L�V�I;ԡF*��9��)�b�OY������'��{X)j.��'���Oc���x��pg����8���An�c�yN��R)��s�Cn�����M��_�i���l����L,rK���k'������du��/��:���;x��{ɻ�o��SOp��u2��{�	Ŵ`�ߣ�f䩧��X�)��x�p���M8�Xs�z2�:d�U��h��ɓ���"@$��*G0V!P������j�l����5���E�MO|��6=�:��}XH�,�^!��C�Mլ����ޟ����-���O����_�ǎR�,Q޺�F�Щ<���QF�"�1��O���+x��%|'����i�ЙN���� A�"��R;r�\�F�KB5cW�X]0�r�cUNVz���DHL,�Mka���B+�ELs�&��A��X��d���~�\����j6`�9B�#^��d#됣�� � �@�zf8FuE9��Cw�{��O<G�\YS�q���i?8�׽��z/���Xq.��]��]�ol�9���*�B�fBV(V�W��3���x���9�f�gX��U�q��YE��r�#�%�~���W){���츂͛7����N�ڜn���c6E��������z?�~�:�0&�p"����A�FO�w4Q/��m��	�h��ғ�NPK�TC���D�L� 1����ٴ��6���߼����YI�c7����є��*����ə����fl=��iI�Fo��q�^f��pks�W�_'YYaz�2�O>�����?�#�>��ϒh���wp#����M���Fc��>�Z�MP:yB]���b&��m��!,:!�o��R�6M���:��Dޡ��h�hQH,LlR���NO�a�r�I���'ף"�n:l�4��Qx&�2�T�\�U�&�S6���?��|���G���s��n�ˤ{{���k5Z^]��B���\��J�4!��++��"�?���6� ��_�y���g�NNX@]���R��o�������+�{�HԵO}������G�������X;���?�Y���
�*��C_qm�E�j�m,s��J�(�%OUC]���4AB���w��e.�~�Z�Q���c��ӄ�Bh�ܢZ�Sq�^VU��-�fE�dVR�X���{���iu	x�ݕM{��I3���jGfS�����C�����'���I~���~�79Q��]kXӆ�^����a�`:.��˂w~��1�6���O�m<�ġ �66X,c��Q��E��t{\�r?���܇�B���!PמZ��2��hL]SIIb�s�JT�\���� �@P��8�-:���B��������|��]���㏓?���fwPI�sg��1XF������>I��}Hj�omґ)���V�n^�������*G��c����i��#?Hu|�k�_�E�昍VW���_B:)��:��n�c�Oq}����b{��Cw�ũw�����R��IMg�׎�3�'��!���ru�+Kh����G��G�d��,�}:IFQ�xm���)n]��l��t�Ͽț�{����V�|�t�崦*���9�g��pŅ�H��]�8�M	A0L��L�wl�-!J0u��1q-
)b�i�����)�iNn3�8}jJ*�
l���<�q�(�\�e�ƌlX���L4�L�SV�!x��h����������;���}����c���7���}�w�%�t�)�#�+�y���6��q��Q�7@��B/��	J���8�)��4i��s��!PՍB����e^wX_�(�0f��b}�hr �3��81|���vJt&�(�w%{;���SP��������;�}�I^��W��먽[�����j�9z�_� ?_;�\P�;k��ud�Yj�j�����{o4�/�z����������4�<#�X��܆�Jy|��z�7��_���3'N�z�����s;׸�����w~GW�rzi����'y������G��3m�3��c�(zI�,A7�e*��e.	����V�2h.�C9�X��4Q���!e]S��: ,@ӿ���U-�*/T<:N��)ˋ�3��Ģ��Gi���xB=�Y�`mݼ�^ּ�7�c?���������b�g8����M
���r��0IJ�[2Ԏ�Ҝ:u���/]}���N���YrIY�Q����ыVՁ�ZN�=�ڱ�<��/P�@���!�/B�ZH�.Y��U1���8E�h���B�G�a%Ay�H�h]ȖB]VT�e�(�w�e�{�����t��j��;�S��$tm�	�+z!0*g���S���6���/᳌]�9{�����/�U�_��R��a�����w7�^b8�q��Y��A.\�����)�H�%_��ʱ��G酻�{���[W��^:�}��\��cT�Vf�iJGi�d�Uʩ�@�`w�!�2�{��댇c�VIL�K0U\L:ˉ�c��˷�qck��ۜ}���|�n����!�p"�nZ�\cK��9
�4��1Q�V)�o<uf(�G'��d�)fPW�t�m
e�ѵ=u��~�5)���l������n",:�r�����@��a��{X=>a�WQ�kc�d­zL�������	Ջ/�y�&/]|���G���Ο;�?��_&(����)FSn]����[(bjš�
�R�"�Vk�F�5��K\�̥��Z�HB ��(��:4�tZ����r���(0�F���J>Z7ǎ�D�@��"����&����(fC�r�&�r>��ㇿ�#<|�yn��}���}�0�%՞-_K'�}҅�s�s����j\f`u�"�Lf�����C+���֠7��������ş�<Ǯ,�w�x_�J���o�c�k�g�?�kso����<�
�ο�Ծ����·>�NΞ9ʯ~�|�kOP#6V׸{�>�r���&�n���^�3�{t�$V��:N��c5J͈����	X�L�j2���Q-J�xAr>���QV%E(bk�\p\PDM���ƶ ӄ�І���d�����](ω��x��.��C4�o��.>�η��ïc�g�'��(^��}�k,׎^/�i���pA!�AY�:h�:u���[�%&��}�]��u�p�W(����I�@�`�a<�0)+N�}�7or��+$�m�.�A+M5��F3�I�*����oB��X�քףM�QxbA�Fb�>�T���&T����`��9�~�q�IE�d�S'�b��q�Ա����Yj+�g�*p����y���&uYS�����\��ש58�QIƈ�����o%(�p{H7�p��9֏����st�}���TiJ2�q�˼���s��0��g4����d��QV�&�*�II�4�tJ�����|�IE5��*p��;!�p����qJY�[B{�x����U�����に�.sᥗy��ge}�0�Bͽ>��v���\��w����ד����(��b����u��P�f�:�O���ϼ�Ir��@/P1�_�3��8©�����&��M�	t{��fRN)B���1�c�lعq�/���Kغɻ��{���~�_�/_��w��`�[�oS�jt�lDcj�靲��$� ��a��h�Q�&����ijl�Ec=ϗ759�&,�\�8�*4�q�i�j5�Q��('L!FAP�a1&�N��x�i�8Q��No�x7������?�qv��5n?�u�����V=������k��ZW�\���yB�}k�Z�~���g������̺=�XB��W�]��3���?[�M���v�׷����_0y�g};��aN���|��g�د�&��]�߹��g����/]y���m��bR�y���$����?��l��Ь��P�;�X�$��˺�y�V����ш�W�!�W�ј���E�M����2�둨��d�,�����o�����w��cA�į�s��'�����ј��(CW5�:^ЕG��R������N��
�r�=��=\Д��[^F���j�$�1i����N��=wq��+�|M(��rJ"+B���ls�%/�x��i���"�a��p�
��K���&(���3K�i�L3�5k�6P�e&�cB)�9yEBU�(���Ģ+��{��U�G�ܼz�;ϝ���s\�z����N�*�qhk)�b*s�����I;�P�r�Ӓ���8�W(�٠�dXfS�Y��@1�0�LY]Yar�
cq�Dl%��%;y��ވ��~�Ս�l�)+G�f`�`P֢mJ�@�(
[28}�c{������AȻ]fe���(&��҇��߄��E�b����{�o���Y�P���4�F�����u6N�aw8eT�ltVɲ4j��5���$0ݝ���É3'8~��?�5���t%~6fYL����)i�bk!�`��Y��<��~7c�����ٹ}�����'�������_z�	��c��tW���?dk�~��l¬��`���$�L5��|�ĐwlSS�$b�~���Wդ-�Q��⼉�`��	�OT�57ڣ��f���h�&�8T*�(C�O��2����|'�9���E���(/���g�����ޤ�H/�b����̇��Z��fiF��B�wp"�W���0�aZ�����������?�~7�
��I*#2����n�*�?�ʵ�w��[Z٘�j��'y��5֯\�����|�{��;����?�8��y���~��}7o�dk�:�r���%S�$�h�	�4I��ш+�Lk���J�4^�2j���(�[��j�Q���sf4լ���ACp��c��=�A'�5:�tsD;w�;��?�~����������_�u�/]�n�ވ�'t5�*�� l��b*���ZŁ6�W�P��-6볳;��["3	��8��	I�᫂�5&���d�����RNЮDB )+����9H�B��n�[��-��F�(�j$z����JqLB�T�xB��j�?ɍ�=fe��`�R*��$��k��(������ԙs,=���Fc�:�w�����7����F���v�;�t�����c����IS���r�$10��:M�U�EI��o��l�����ل�Ҁ��K�Z��v��&:M�z}t��[!Z����p���#�����Iӌ}W�5�1���cw�-�s��ȼ`4���Er]m�\���,���s�`*18��--�]�`4ݤ��J�u�|4d����pl}���m\Yr��y�~�k�,E)Og�C�gl����)I��y�!���&ϝ`�(EJ��:Ӥ݌K��[ܸr�7|��|����^�g?�e�y�"3��WVY�l"��v)���>�4��T�GB���XO������u4�:�0�֍���L�>O�7���E�j���`��Y	jA<�ֈ���V�^o���9{����w�oz_r���Ǿ����N���eg<�!˯�z�']��p�sި�M�Z�R�"�q!�3��/��^��@����?�ٟ���?C�%�I3�F=��0T���[�#+������;;��k5�����}��/q����^���=��?�?�g��W.q�{8w�<�k��7���c<S�rV�@f���W�%��+�Z
\4>�	}5_4�b��6�Ra��h��c��RMKʼ�E5�&M�7�r�wEIQ9���t�#h�7��j��w��#|o}�Ä����_��g���Q��Y�M�0��ylY�E�y�6�5��읣���d̪�F#9�ɔi�uiޡ���t��ޓ%)is��wk�ET�R�����J�1n8bz}��(R�1Γ�Џ���V���y��Ʋ��[M�p������I�]��$	^k�Q�$��%�&��!��ɳh����RVI��}����ࢢ�1��������$��)�-BY��<æ����uA��Jj-R�P��(1:���u��
��P;T��m¤(*IH:9ʚ�U1<�'9F[
_�_��POY�$&a6�RLf�"�&H���MhX����� �.!��)IIݬC�7��W�`���	�0��mC`\��UE��%`�A�hC����fXk��I�G)�xn)������hHWC����I*O�̕:��Ja�Ƙ�-1Њu�[/]�s��?��c����#���}�7�r��}��|��+�唼�%M,Kk�T�c<�����t:���"��Y��4���\�ع1_�6޵4�ŢU�����I�*vy4�ZEuH�*�W��:A�9Y'g����fy��[������r���g����}���ϑ��Vy\0\-f�O���+�?,j��+�����)C�U�a�v���m���Dk���_�[�7?�S��d�O=������⋥��u��^������ݱ���q����ӗos�mo�����{��&^������׾�4{�[d�X?��#�ʊ�����!�񌽝=��F�]7��J9
\�
J�E!����K�!�$6��`�&���G|*!��u�/� ��4K误P����,�������|�������>�>��\��g�7�K��ӢQ�R��M�ƇX a�r�d���kj�(����άàÄ�t6������+���c���̒��I1�*g��ct$@�XR��ј��MқCN�9���ړ�Y�S"͘H�1�F=4ަ}��14�����h�1s��L�T�Q���&�#G�,�i7#M,��X�1X0�N��ʀ�۷pΡ%�(M1QO�H]��q5e�5���8�$��5�[l�ı���ڣ�n�O@�����̐�R^y��rF�e�tgU9D*:ڐ��B4vZ#�����q9!Hݔ�U�4%�x����R{n]��h:�XC]Tӂ%7)��ӳ�ӈ�8D�f�E�k1UMS琥$�>~k�Nڥ�K��y��K�[{��EE���"�����g�^� 4����K`��/<E�c����/FU:��+�[[ȭ[�u{tר��=�b$�0�Py��^����ո�|ZpD��}�}�|���>�0o���r��A�{�_z�q�z�i
[�l��t�d��ɔY9���Op5��[�͢�MU��Y<�ڕ��a�X���=�&PM�kt T��$��A0h,I4�h�)��!t��(g��x�������8���e����d牧�o��t�FLnNf#�:�t�g��QU����ҡD3�R$9u������[c�Z�������_~���$�<#�p�j�Q�
J.��Czt��qY���i�m�m�v���^����O���'8��7���G��w;�x۷��s����1ܺ�lV�e	�6X?~�,��17o�dow���(���<:�C\f�)�{�ܢ���*$���YS ���y��ji��LeX�8��5E4�h��<!K��P��.'Ϝ�]�{�G���<��v����/p�_��t��Y��d���s���%��0Q*����` ��s�S�*�i��;[���;q�׹���\�q�g�����{�{ｏ��J)*qL�3�x시>�$�<�/ӕ@�<=zZ�v���>`fST��lSs��&�>GT#�s�fK`^,$��%`�!�~V�*���6~k���/߸̅�������7��{�k��t�v�*O?�$GΟ t���2k�;]�h������E�fs�Z���Ӝ�����)��!_��gx4�9{�y~��?�w�^��J�G����)�|�G����x�k�q�ߧ?�(wwٻq��n���I$VS�f��}n}�q��z�.Լr��N��+���MΟ9G/�1^����S���ן��?�}���&��tB`դ�^�J��͆Ip�I\�5���1i�7����J�|]�G��`@9��+�r�q�����_����$/Iz���&�����������'H�9��1-'<�;_䉯?�G~��7_�ĲM8� �vo�ҫ�4�ܴ�/��:M�	l��-'；c��cg����W�h��W�Oj�sQZ��;�>ͯ?�,���۹��o����^�z�9�}�;{{�1,�Y[?�'�M&c��!�l����>
QlJ)0��J�E{��ĢT����D�M�Ejs�6���h�sQS��6���=B���Q8�đUy����[����o\��O���שw7��1}�a{ݰ9�N0��cG~���^���kc�lB�w)��nN%�������u��3�kD����O��N���&�2(JҺF�ό����w����7!]���i]��=��N�뭜z�[�9�����K<��lm�rk{��7���tH�9EY2Nb����l1ԡ(�E�Z�K�f�녾�Aj�r�%ԎZb/��StjAC��tzZB]�]�s5
8v����7��w�����Ey{��_y��>����[d�#V�gM��՘���-�aW݄��<5��>�����E0C������ʓՄ�������>�̧)|�`c�������ֲ��F�jF�1�w�Y;�����H5���|��wt}��(7��;{v'��d�#�B_[�:!&8�=:�٧��E�=�ЛaQ���!�ɖ����e��RH`�Y���&<t�O?�U�Z�7�w��_�U�;}2e蚔��m�^���>�#�z��.7�_a-���c���:�g.п=䄷tʀ�Y�n5e��*o���2ש����ԕG�����}���3|��Cp�P�LF#:Y»���>|�����,������s/�^���hFoZ�9HM�W)���٣�����<}�vww؛�yۻ�E)§~���"�0��{�N������>�c������ݟp�㿅����̑�f��g)����a��o��>��^���[5?NMX8Ә^��p��pB>XfǗ�ǉG ��;�ů������<��wQ9᳟���[���6o���w��3w���'�g�W%�&�x�e�'/pjȧ�ո�0Ɛ��'	[Vq����}�{|�j9����]������fl��~!d^3�	��+~�=}����9��w���΍ј_��<��ܼI)�`Y/'�d�`:3�L�9|YRLg�N#̽n0:aVe�(��CS�¦�����*W��Pɒ�nڡcc$РPX*�t]�ז9z|����u��7q��*��=��/���x
�6��됮�II9+��+��O��+U��Q�Z#��Yb):�����Q��/����+��?Z����_��o�����G:+�ޓ��A���}Y~����,��#Y7C	��`��I�cp�9�<pg_�0fu���m�o�q���x��<�e�^��!���Psŧ����&��t�Ǽ�6�\�C\`)�j�GP�i���v%�U$�"� �q��QN�8�����{8��s�K�~�9v�{���u:�)�ʑ5�,�uM� 5�<�PM�MS����Alh</O*����5���ű��.����+�>ɳ�>Ϡ��׿���._{�	�ݼNUW�4���Ӽ���LY����s�T5jw���&ns�tV�R8z��t���~�a���)�E1��c!C��
����yDq����+nܾְ�*�w��;~��\�y��]z�lc��?�(�[;����5|QʒzVr߽����������<���*յ�\����ئ�=ᤤ�I(�5H'�y?�؏?���<��/�?���������\�p�[7na-±�5�;�,�*N�[.w�\���dFwg�A�ȼ�U�z�ˆ����s�W.�Ȱ��殇dwo�O}�����$S�~��>̱s��.��M��J¹΀��k\���ȷ�,W�����g�� �+cn�u#��Z��AM���`��v�P��3&���)�w�Ü<έ*P&��yK'O�{�'{�_�:F+z�.�Ξ����fog��p��,�����_�L��6�$#-�8K\\�>'a�������� 7�x���B/!��ы�)��彂�QM2��.Pja�)v3a�xv��l���7��{��V��>��Ɉ�W�r��U�y�%�ܺ�p:���us���F������]-�d5�%h��8�T�T�5��b>�TLɉ !`�&�	�2�:�� (��.�q�����]<���<t��t\��^d���ؽ��KWX�:V�Fꊡ��^�n)���6�/�����o�JS��(&�.�R�E���[t���Kk���/�ԏ��32��3���@���6�ݱԇ�������������\�L�T��tX��'x�s�=@��;qY����v��x�%�ܸ��h̍۷�u�&���uB��b"Jk���Ԓe9(��]3�MJ^p⩽'�Qz���68ut�{Ο�̙Sl=��R���6�_���g�a���KV��lR��̃����!���nb����F�+W�ȱ�ޘ�.�^ҧ�e�x�kx���	z�Ó_}�K/��՚N���U��C*W�����@��૊T�Hށ�}��f{�l2�Sy��#�(',�zt��V�ΟZ�b&@����ņ(�G�}T�p���x_ny�o�c����ԅg�YL��+�7ֹ|���! �1�9{���U�����X���I���O?��$��,zRal��;��U.VS�����	����[ń��`��g�R(��C�g�K]�����m��F�+7��بj��}�.��	�q�����saB���M?�Cܼ��(n��0	��l��R�%�<�IY[ZaZLɗ;���@�MH�����Ӥ�{&5y����&�
�h9TP�����Ag�Ǽ�н�Y��x��WtWzL�d���q��p��n��{��:��?�1��c��m��e4i'!�zY�r�vG�_����&��}:7v8I���fto�7�5��r�gx���i����?�I�R�4��"ߛҹ����	W����:�a7�rK=�0���7���-�p��8��7p�C��Vٞ��~�*.��KW^���mF�	u�X�nM; ���&��m����{OQ̘S����r5�ٔ�(�u�v�A�qr���q'w�y���ǏeE���u�]x�[�}���+��!�T���x�R#�7O;~�P�c��Z�2`�a����R���FJ����_�������5������%��gtg�ʓ����D�y�xQ�Mf���/Y�䉸ZMql�
��Q��6{y3��wRg)��xW1��y�&��r��׮1+J��1EQ1+�:�Z5&���UMU�c��.ݼ��	Y�1X�s��q�:s��Ǐ1XY"ъ\��mn<�W_z����ݸ�LF,k��0UŊ��.`����[sBP����(Q�-4!�n�-rZ�j$ u��Lk�+Kj�l֞띄��1���|�d���K��y�Zf�pu�xOoi��h��%���S�ޥ7��f�{c�QA���c\�jM�w�Ƃ��&J�5ȁAױ��4��i��4A+*L�C�����;�;t�����f=����s�Y�\�ȴc�8������IQ��Љfiy�e��GT{C��f{�loBo�`\��9)6��-�v٦fS9V};.�ܘ�u6�13q���*
�:]2�ɭ%њCuk����S:�1��e� �)N4eH�t�&5;�s�ͯ���ތ����m��2ǰ����v;�wx��M��~:v.\d���X�x��m�iE�+zƐ��i��+�kA�����:@Pz�
�b;�e�p�G�� R�W���%��#t�=f���f悔cw�G<65�9s���Ĳ��%^���t��F���wY��j��D
�l��'�p�Y^��9���|��R��d�j�c6cm&/\��t�ި$/x�N-U�0�3q�4�&T�2VB���O�b垻8u߽9s}d�iU�}����\�|�[��L'S��1E3l)(�*��J��utS4K���&_���&�\���cGy�}p��;�,/�Q��F7n�s�
�^|�����]�b���ᴔ�S�J���KO���˲�~ۉ�6jTJ�)��4	�ۣH3J`V���_��o����A�7���?Nb&x�dFg\�)�� J�1��*��U�G���-=����Nޱ��F�Q�K`�4��28}�����8}�����?��w!1�^��$PU��,(������jG�XkI���U:Y��I���*d4ƏG�n����|�%�7o�GCR�Y.�~�RcT�	&�$�ޤ
�4ZR��0*��uD��1݄��Lk�$�t�wU*PkO�
�tFB�.Q�a�4��.��
w=�z������L���5��d6�������,��7�?��J���qI��r��j�n�h�w��
�A��Q=0袢A�"1�b�����%I�n�Sp��E������`c	9��V�Oap�$ݣGPݔIY0�M�c\�,�
u}�rs&3������"`�5��KUb�iM)�<��-g���_�AΦ�������ʂPׄ�B�3��:��T${fwĠ��U%��ȴ�\@LJ�&5�4�±SY���Y?a�)��S<��%��锕��ј��姞��NIw��;c��)�ʒ�� �ȭ�]���!z��5z#��]�^H��
��ޕ��$xlf�9����w�G�?�����Y�u3��y��K��1��Q��O� �ɵ��~�E�q�ޛ����%+X|U��I�c����R5������wl�/��2�d�&���H�d�ы��[;tF5KΒyMY�q��eh��j�G�&�iƾ��'�}��&�|}���'8~�'Ν�w�8�A�}��mn��1�ٔ����ۧ(
ʪĹ8�AiE��,��Xk�t;�,�Y[^���`��
a<�������l^����&{ϿĒ�d�Y1�\�0+��N�i��]�m�Z�oTN������U��b��81̲�"�Pk��s��}k.��h����?��Q�9�IA2+�}���^0�[y;���Y�ƎN��Y���ʹ�*����`:�Y�Koe�գG�Gר�;t��Y�X'_^�d�ƤYL�;�OM�\M���ј����;���ooS��Q��g��*E&�S�t��{�Ղ�S��qb�w��1b0�h�(o	�B{�U�v��o�fo���u��&P�@��[i�1Y��L҄q���%�'7����r�Nb]����d�ԁ�N�U����t��D��h,TbH���fҝ��`��ӡ$4C?bs�Y�,<DMP�@KP
��uع}��DCe�b���r�S�){�}H6�謭RC%����kz〽�OZ� ̶v�z��[:/$&��=�ۉs�C �R�g��:tOc��^]¥��r�N�j����N+�I��d�q	�iU3�)ft󌢬p�Iht�P�
���jJ��Bvl���*3+t7V�-�x���N(��Fg�II2�У�5��creȒ��X�|���H�6�i����ֶy�t1���FaSK���T%y�Ri�8��M9�a���_�:�����&T�)|�h4B�@�3D�K�"��0.�����M������B�mʎT\rν��~�-ܾq�N'���˔�I��*���#;��S��:�ZHMh�ȟ`���֔6af��2��"���0���$�sz����O�=�ڑ��9Bwu����t:�,J��F��Qڂx|]�
����ߧ�١���d���xk��pW�HUa=l�K�I��������W��iR�����^���:x�A�DSd�Q�0M�(fe���+����x��5��������34B�=�t���N�| �A%!Xdɢ�V�os^�V"ߦ�tGB�+�t�`�G|���Sal��xIj�;�8Yi��mm:���U��P;|]A�0>�������Ȕ&A�j��5�+�E�u���2�1$Xe���]��FD2�W M%>D�ԦҶ������\�M�c3Eb��)M�j�ٯ��>����@L���0AH�'q�?�5AHc��\��~-Q�x!�&�����|���p�%Y�q>ԡ��w3A����VQ���L13����A��P3+
�Q��8`kh�Q>��`CT��r��[V��^)����ɠ�"yJ�����c|�7�ѝ�:
�(����X�X��g�F�󑀷2y�O�����Hb��ǅ�0�vF�IA��1k��ǻ��=� P�=S+���H�&����fށ�4�Vc9D�_��r�z��ÈPL��!2�^���cA�� lV�F3��#�I�q�H���}5?���U쇊���S�8r�.��M�W#��LP�)Lf�ʑxH�#�	J�5�^k*e(�����Z��b���)�&�qb�Z�mB����$�.&IA�f�SAkl��	EE��PeE�R�(�Ď�!xO�N��@�u�W�ǔ��z_?$�8(k��t#��&��C��LU8T{���omx�ߔ֠�[�?�����h �t:�N
�ʑy!H�Er-W�CZ�[��Q���h	R�7�(e,6�Ȓ�Lk\U�|T���S�QPB�X�Gtk���Q��6�֒ꨜf}��@*��C{�i�Q���/@�rQ�C<����`���r���%`T44ZhDr8�6ת�H�&HҎ�n���G�T*%�V��$if��fh�`�`�����6�� ����ɽ�\��b�����}����^�_���~\�+���VP�(U Y������*��T �X����¢U�p�ܼa .�A�BO��$����4��^�kUZ�l\�%*���i*��xp L�ĉ\Dz��k���
�Zt�R���n�rYc*�{�3��fT��s5��5���V�B<��Sc��
g�+��Ŏ4gS|�n{FA�FF�A�	X�7�U5�r1BR	�l��#s������y��Ǻ�'t���<��6B�k�t��L�e�L�����Z碆�1�I����BQ�i&�F�Pᒔ�jj�B.~���-���4CV4Ts��4Mc-��������Zj��I����:���s5�X���SA�h�7�Jk*�0K&I��ZJ�k������w��-��i��!?�~���ړ�*�ړ���5A��	}���.ϛN��ޡ���Y���Z�̪^�7�Q�Q�jc��JE%'�(%W�����c�=�!��DE5�T��6��E�k��DF�u0�8O,��ޖ	�i\�"UT=G���X"�$�m�s��h($�b{����p%��R
�Αt:H�H=o��Ek�j�lh2��5-�Y�e�%����W�%d��W4�2�C]�BK��$�� �x$�Z�A5�
�I���ƨ�8����ܢb!�G�+�҈�i�@4�B�3bkaR�o����yH�$��ڂ�:�ua�8�
*	��ū�q�@"��sh5�6?c���U�Z+�Z��ׇ:	e�/�ah]��^�Ύ�Y�K4�y�c����ޔF���J�!o�鎠���x��}�A�C�vs��Yp�PiJ0MT��wH]��:
?I�8�8(�6�64]cc�J�Z�҈MbZM)<�ċ��NjbI�V���iDiL�Q9Ođ�*:�\%AŢQ�|c������0�����7V�P_����3QO�Iv�+sӣ�A)�D��(s&F��P%	�)�s~�5�'��������:Y���u!*�U����e��6�C�����HW��F��F��ir"hs���T��q>�&H31��Zy�������	AY�R�Yktb�����:�<��dʤ�҉F4&h�D��5�nj����A�>�gJJ�I��t�%/��?�6�ׁY=�ؚ47耰��v������Mcx�����ԥY ��sC@��fjW�$Q9��J��"!Z\��9l�y��Y�jI]P��������@E�Z�8�}n||h|�C���!������)?��*�_5�'��U31k�Y�<��5�ه4�{��T���f2��(#�a���q�����R:��&.����V2�k��1.N��h�~�F\�6۵�`��=T<N2_0�z�����i<���<�xα�4��8(��>_|)�KL)��V��c~�(rc�C+@>DeGњZ��DlւM�l�H�B�U]�ʙUz��uK��.H��d5ʠ�V^)%Z+1F���Ji�|�����Z��Ej�OUm���Ė�6��bv_?W0j_�Y�f�qN�P+#�2��RhE��Q��0��9/|��6��{Jkп��?~�A��Α9G���XJ���xѓE�Q)��jH1A�M�\����Cb�ee$����6!h3�kF�u�ZUZ/+�:²��zW���\�,�L�c�R��,w��A���Rk��+0�pK�%jV���z8E5�@�5V�P+�f�.�h\�0[FU1�\�bӄ��Ja�m���Pj;'	QB��&��O�����b���k�o� ��Z���b���!C�b`����iv�5�Xֽ0�1���C����s�UAU/���m�27\q50_�D'��b(t�QdDV����nB��-�D#�o�O!9�o�z5��c-ŁА��E�c����Z����f��E��<�/��\�]7�y$F�y������k��A	�P$h��V��!jq3���9�y:d����J��ij�dF�jq��ڗ*8l����8k)��6��k(҄=�j4���FWt�o�����^R.�D��D� *&O�ٞ/:(���:(<U5]("�|�
(�P��E��ip@sOMT)4igt����4���L���C�Z/����ƿe��������C�sv�	�+Lq�S�oף\@�������Eo���J�pTSģBE�hK|?���T���B�1�`�|�谪�l����sd�]��ο#��8��Y�xA�y�P�0�(�wٺx��ސ$@*��4/��b\D�w/�90^�$>C#��k�vsIYY���Պal�1�v_!z���N�1�u]��ؾ���{|�\2V�&���TK�ۆ�u΋��Z�!^+�1��� sϲ��hv�7���oE#��q�5ˁ���Q7�G��p9`���1�
b�D#&|����,mi��|���A���(4����)������EMT@�9�Q:;d�U��<��X�h�ۉř�(͒.��E(Ӵ��,���i��X���o���h
_c�9kg��=~�]|7'�)^�dkk����K��F�
����V�LD�LP����8O�䃸�|RZhBA�f	9��}$��j������,�������a̌ƛ�x�EU���'h�������K?�Q�4��7:�'=0�V��x�0! M�y�Q(BBX��\Ue~�i�¾iŒC�̍@�Zbj@�`8��Z�J�F�45�47obm��w�֞�*�
(kzy��G�ck�+�_`���SW�M4j��nz\�tA�>�hMb���%�p�ah���R��A��M�����9E�h�;d��з�"_�M�ϕ���Y�SŉS� F;6�$4�%���gXTi'��a�0nzqQU��x��1��-��/^�(P�l�f���Nk�4%�@��8+>ngc����������.M=F��ik�%Ѡ��D �X����r� k�áEY͚Ē$	����5��[�%����i�ł0碈Jpq�ԡŊ��V87�֦1���I!�m!D/�+����J���m ^�1�Pe�P:���&���[E��
��25v�����]��sF!�9�@��%��/����q�O��ߜ�/���b��!u��xU��<v�pZt-,�k�����V7�(��c�f�P;%��ͬ���C@(k���k���^�Z~�i����O�#�=�R ��,<#����*��a��d��kb����;��s�=:x��x%d���d�<K3{Tk������?���L�m��u���j0J��ή�l��P%���PZ�����U��CQ�F�:�u��ڋ��H�%b�i�UP*�}H}p��B)����t�)7�xZ�%�T�JK�}ڋ���Eš�Z7�H8���y����<>0��T�ؼ
����JE-�Mt�e0Z5��M뜠��Tup�ѳA#Fk���4Jk�T|S<�{	�Z�n�ֽ,)�H�W�b֯���AB\;���V���Ҭ)E-2�'���P�a����J�U��s/��&��UP(���C�h��I�̽ÀR!�ص�jJ%Ɗ1Z��'x���'A�5&�N�sdi*I�JQV:*���Ō*f�U<�͹/�H�:fݕǏ�h-��Zlb���;D���Z�h��Qh��d���n�:B��hl�6���Q_��*-Z�$�V�*��AX?w�峧��R�׮�����c��k��#�էk/{EU�hV0)+J���J�`��V�w�w8t����#a���V'(q�s����KY˷�֠�!�?����$6zVp�͍��+�	B/�,�:t��4!�J[��Bf�4E'�T�|(k/E�BQ�zV��R����M��(!4a]�����l �� �C�y+��GP���˺��h@n�?M�2͛4����51�y�����+Y���?�	 �q�l\=��Q�F�a�9W�P�pFڌ9
Si�^Fy�����t�n��<�C�u�l�i=������w���?]=�r~X��N������+A�$aleS��A:^#�ѱv����}��������Y�������t��纙4I�X�#�2p�0����l���?lXof��|Vo�b鳺����Vw��x�>��u'Bӷ\�H������ft)*q���'KSb�����yCD�����O�Յ_�?����.����3�kD�*���a�q~LP}��>������2�)\�`��;x�L���a��d[=��	+xwe�]�����Y��8l��&��i-Ř!��^�����=�0m*�=�%-�a�]M�����Txx�4��%�B'�pXw�<�e{��BIE'|,��	�غ�)���ڐzqJF9��{
��6D3j��C[y�収���(�{H��
L����ŁR����[4R[@��&�H�z���flne�6�r`5ݍ��Qc�n�����:m@�LtA���Es2��r�v�f��OK��ȄZ%�LA���,��k�+�`��sPF�SO�`H)ŗ5��8˧JU6o���n]��{{���'	o�	'h�o�<��u�T�g��f�ZՎB�����{�H��]Cĩ�y�	�S�;�4shb��C3�8��:��`��'s��zv%~�cIO�}j�&�X��s�Y6���M
���U�K����H�vr��J*
�PZ�)+�M�|�B�/*�-"����bv��	%��]�mN�L�u ��h�eho�g�`��g����#�&�ʮM9�fw��;��9��M:��K,��>ѓ^.6�1��կ����������w�خ.�A]g�7�rD@<��&C�D��ZvZ�ɜ�+U��}�!��D[�W2�W>إ�&J�8���nk�cꖷ���b<>���H�k�A�=�)�z�u�Ke}�<��
����Y'DG�Q�ų��#��k�+)W#�'���B W�Ҭy��x��]Tw��s��T����EM��f�r�����7�ʖ��h2����^h��S��ly�N�U8-t�.�Q� p^���Zj��
��|X�{*٨T�$GG�����]�^�7<@X��$������CKw�S[�Fb��ꬄW�Y���}5��"Ū�_,���VS/P7��
��0���*�=����+*�h0E,[j~~[�����Ie���Lg,��L���"�?��O��� PK   ��X����	  P  /   images/471995ad-a105-47c5-9945-45370623043a.png�VWTeai�R���	EE��Pŀ@��P jiF�J�J@�MjB��B@:����Ĉ˜=���7g?������y���n*"���17����!X����t�qfN!||
���/o|�l��xcG�-�O@����o�_�'����X >>�ys��]X�z�-9�lI޴k��5��v�T����L�T�>{V��6���褠��.��cG����aP�]B���8(M�L0��s���@�Bݔ.�tQ��po�W��_����A��ނ<�5.oxW�1T �ӸӮ������Vi_=� �8G%����4�"�c��(�E��^G����"[�#"���K{�k�֧W��#&CUr�E�����޽�X������\�R�8�<ui��m���g?yg�N��[�4I�g�766V���w�I4ՓB�"ٴ�ȭR��(7ooo/U�����H}m�FM]�jE]�<EEZ�-ӳ?żg,��!�@�̕��e�8���brI�^��|.���Gs�j�Zε�ow�����0�l:�l�cCB�^��\i��}YZ*��.��dlBoRj�)�L��_$��{츑I@.QC�b���>�1��ũ��{B'��'�n�|�����+=�v��U�60�M�y0�M�Y0�4u+xa��T��U���>��<����	�4vw=]|���%պ�;����}����o�em{�J�Vab4�����F%�f�Ɏt82�i�e@ �P���Eʐ��l��������èV�M���\c��$uI���?�;����˗��+�se��Y� (�� ��e��<vr�/#����۬h�Dǿ��4�z�Yx�Kr�'`���z.�Xb��4�\&8����?�g�^��j�*��@'��%��l �����r?�}��[p>���_5���2^9�G�VQ?Ӗ�� ���:_��?���eoՅ>$��gըOe�	H3q��9��G�?�E\B.%�m���D��K����r��k����e-�b���)���m]�Jǩ;C���ӘM[>�o��[�Yq��#m��ʏ�B�G��>v�gB5��?i��&<���������R��G(���l�eU��i�$�����Ɣ�|�W��H�c]�Y�^ubU�6C�eٌ��������Gs1Vަ)��e�`_(t���"n}�����@�;Z{*�C"���P���v��H��sC��E�R�����q�5��ee
`���^��j��C0���H�́���_�{:������i �ɱZ�}�ibZ/�3!-���b�n�!K=�V����I�h���BG�#@����	?֒���Vl���t��-3[�?�.z;�[1ѽ&��]t��J�_�7 '�&��}�X���;2%�|�D�ӭm�;y��U�<{�+T^ZW��A�]<�剠�B����dxs�5���I�J+�#�u�>��]�^NoeM�^c��(�(�2���a���{'M/���{�ɚ�$�KN���5�W���v_|NH����ZV�,����\���0�(jA*©�)���8 �1�~R��j�����x�P���{#Vm�>@�\q�Z�\�mU��N�~
t���c�VL�������q�a�9��4Sn��`%�% )���]H��Ly������	>e��G�O�/DҤDL����7�}E*�l7�t6=�uJ=pO΢U�(Ɩ;�@tsM&ہK훬wOU�y;����f�%������k\���	 O�n6dBth���3�Q֜�+��#�� ��A:�~�~A�<u�
'�R�(�i7s4���VM�$��;��݌�;ȭ/������ȩ�"�
��b�w-l��In=jՌ侉ڡ��ED��G{,�-��O�ɻ�0�l���%�˗c��+׵ًm�Q{A�5B����u5�ͧg$�#���j��!b�?6Kq���J��3т�����m�8�<"���>��N��$��d߶�;��7$"N����;]x�It��\c�Q����m��h�z_�f����2�:��ԍ夰�����عH���U�m���h��V���W�����������&t�,�=C[y��^�$!2���������u��EVs����ᮘp�Qղ� (c���U��7a��*�����'����{9�h+��n�x�ۈ_������əwg̿���(���9��?�V�L�$���A�w/��Ƕ���~IN�?Q�?}��[K�����ދ�Ĥ�Y��lg�
�� ǂC|#c05����:ͫ�Ɲ��_�%8Y��Jyv��%�-n����j�e��ؘ��S�!M}^�N�j?�G��Uj���}l���XOZ;�;g_�FL��Y�-0s�#�[��Θu�<"�wv�f�
|BS�wy.l�[g �l�/������VM��iU��ٍ�m~��?]����׋�gn��A���PK   㫦X����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   
��X���Ʊ N� /   images/8eec4e94-481e-4d4e-9432-645515506382.png�{�S���6-���C�8,Nq�"ŝ����ݡX)^��n��w�����S>����=3��d�;�ɹ��I�?��b������a��I�����|]P��m[X���Bu��u��c�}]�x��y�����K�kz�v!�}��B�g���.�>�P�P��^F��bn��NgbA��AA�D|��F	���ě>k����|�a�P�Z���-P 	�����`hx�?_Ez�����/�ż�$�?����ڢרG,B1S�O8��ۑ0���5�?�I���p1S����_���vo����/�L�����z�XA���x��b�o�ǧ�������ۓ��ڋ~�F�����b��r�E���T�0�k�>��:"�y�DR\|�����{{
{)��`)�>�!-�r��Y�mG\Z��t����	_~��a�.p�!��4�y�VX��Ǽ���Ï�K�W��GY8�:��3�%vWpҫ�)&�z���#2�s@��iH�m�y�G���	��{y!a��-��vU�l�Tajй0�W�vs�	n�m� f~���S�qf�8fƪ�]C���&$�;S�O�y8͝��Ȓ���-�-���Zʺ��5է�p����@�i�ɓ����cQ��7ܐ�Q1�;�&��Yy�<zΕf;+�=�(��r6'F�D�tT����
���ÅH�V\� �Z��A�Gt@m[��#�-�����ޕ&���[�d�9떝��l�C%1�l��&9�����}�CU�BO��}�?����_��s�:�eQ,�:y��N32�3%���ĕ"�-G�e;��M�CV�u���zɱf�G��|�'�a=�87'm3��� }��\Y�I�=NKn� �T\Ot^���P<�L�~��r)Wl��L��>qO�V�䦉���s����]�6��Q�j�Iǻa�&���*�8���u2�/!�`����KG�X��O��<���]Z-;���Ȕ}�ann��bڂidՑ 3
}o������d1Y�|�9%u�5{�Ϟn���`�O��T��GW��,��:��6�2-� �VZ`�1a��r(�z�ʎ�����D�@�b3� ��ơ7����e�Z�
� ��A�E/"�p���=͈P��d-�)��%�T̯��!D��Ϸ*��  �?�%��a���3G�ք#���I 5�R��)�;���R��f���kjta���t�h-:Ek{9�ۻ����ރ1�f0��*mO����`���d ���Ŵ�����.�g���?8�b �;��?���Q��ìH�B�p��S�IH�c��F�W*O�7����g~����>���1�^�b�c*+5�����(&/M Ֆ���74�Ŕ�jD(�ĸ��UP�bk��/�&X�7�u�GBa<���;/��� ���DBFt5G����
�"Lb~)ѓ^��|��=%�iOwp��6�����祾.�yn��b��ێ�Wک���>!l2`�T���+2b���g����|(��k*�J�%�~Dm~No]0,�Ӟ�:[���@���2��{R�+j8�,��8'�3[��{YR�|��
7�2�a4$~scV�h�F6��.3A��U�=f��i�o{��P��SB�!U�D��C���})��MGOO�D��&$_ss���PX\Tt�	��
/���d~`�����i�i,Ҫ��o��:������6���vf�e� 8����q�P�F�R�@�SW��b��.�y�0�Qa�I����a��n��6©���J� J�x��zp��5>[�O]KCC}H��*NeK��C�!Ry���S4+SϠ�~���1Oɮ��,�n{qF�De��0R�����-�|z�s�?�:��G&	g��������Q��D뾢!!�D���k�i� Dɲ�6~w�#ٞE�ĭ������0��iY4Kξ+~�]��-EӗH>�=*-�3�y;�4�t������a1U�^F��ܺ�gN�]�a��Q%����HK��_����V�[a�a����a���X���ŻfNv��fϦ)ۑ��bUB��e�B7�dW�?5�~�[R�kh4{Y\��|���W��_����[�Ǟ�i�cc�Y�R��BIx���:�Z��5r����'�����θW�(X���c_�ٽ+pjހ�����SQj�ڀ1Xy4wr,�!�~��s��[�;6'���.{�
�|tK	�P�a�G]���3��SJת���������5���n�1�(�A��aY��G��'a$��<ӓ7��DY�u{������n��r�էR6Xq��iզ��Ao /��$�6�������W>���y�	�cPO��eP�t� b�9��B5+5��5}K,SK�c̫YmA�g�:�7o�x|������&��>\�
�0�ce��8#h1���H�|�tw0s��y3`�p>��~�x嚋�9����zʎ���1)$�Na���d��g��;�D�{�o��wS�v���p�%_��}��w�&y5�-�q鲅H�~����S�`�P!O�ȟ솓�]�����n���qu���\Z}�\3�s��1y�)��_0(�
��1�N��d�c�4�k�R�*mﻈ�3h:R����L�/az��t\��l����oV��+
��*큼��Hu��)޿��4�f�QI���<H�Tk*���mﱠtJ�O�h6�銘�Fg���.���k�i��dG������SJ��De��89x"m����T�_�q��\3��C��+ÿ��v�[%��F���=�@z{Oe�Os���f�7�|k*|t�-��D�U*������6���N�{�:7�!Z��
pD}��~�
���߲�����ל�9<s}��ɚ�C5Ǔ{{�V7�Y+]XyO�O(���(F	p2����Wi2L�ȳ^B
:ƃ@����o��(�w���W��d����FDVZ�[��Ca�U��5R��N�n}j	F����Q���X���N�Q�T7+���9�)��	!�����ُ�?w�y����{g��Mvګ8��'�s2���m|�<��29��˓���}ʷ������*����j���������N�6ͱ�w�C$M�@���ӵ�(}�Fj�x�
P�`"3��t��DRI��c�4N�QkF�E����[tg���H���+�M�)�+P�����������]5���n���HAHO��z�<�C�UZ*tc�TJk'��9E0f�`�L�o1Ґ988�g4�@����"'K�T�n��΄��e9�8�ݺ�g>|�A6T��2}J�5'��d��� ��_�{,�vMۦk��kF��G�h��p
74��x�片�x����W�c�?/��~gS+�h_%Y����N�3��mm�E<,d0�3�D�D4F@TS�u��P���#�t`���V��D�X0�/yC��{rJy9g�?������#k��n��l<�'�7�cdQ[���mF�e`A��^g�|~�8�*����fr�v�0�]#��f_6�@#��
������������?��[b��G��ڏ�Gs:zƒ�Mn+CQ��ӟ�L����P��e��39��;�D�.�N@�n��h�h�"s��d0�D��Wi��
�b~.|�Y7~<g��i�jG��ǋ��O�H^�69H�Asnt(�Ho�=���Ǉe�����bSc�)�n��U��W_��8�8C���jҦ�����hXo�E��EzJ�ܦ�#��S���&�B]a � ���H��8��$:�I���r.�~��0քiy\�˙n�K�@���mF@�ڥl�=^x6�]�3G~�}�FX ���P��$��l$G�?n$�!~�Jfe8sa}FLF��v}���@���]�Ԧ�װ�?!s�����'_\�����O��QzJ�Y�WO.عl�m��+�>��{b�ש>߼v���A�W]k���'%�L%:�$�'غ��嶎W
���*�y�6�7:�HȐU����%O��I�.�Y�Tiv�|���rl� ��2���#B�{���T����i,JvZ����|�
ƕe�4C�y�+��!JvǢ���!�jһ��c�1���	v�1���ADtjk	PC�4'�׹� R5�O-D�����VΰPci����:�02��7����%^]�%�Hh�Mp�MG��d<m��>"b@ݺ�&�N{���SbT�q[(1�kȉ7MK��U�����[9�|���$����~�4�୰�����H�C*�ۿU�'�P�H H�[�(b�����/�<FC�[;�$gJ������s����n1��/���\4����:p��bo��~I'#�v�`�1��kt]E��²Bp�6�J�������/sr��,��]T�;�~�������a>B��炵m�d}�����R�vy��8x%�i�QLdl3�Q�|��X�'��0����~i�I�"����q'��=��B	?��;�b�R�e���	אּ�]�6�)�pG��/�LR,��>�8���"�_��8��)de�.�'��?*���;��z����\ȫ��̄V���0�|��IG+0֗����P��u��HǠ��>Q��ͨ�=exq\��M�Y�`F��$�:�d�r�<��cף\D�5M�t]7����CHꢛC���}��b23�Yt��v�JO�K���O�ғ@��+o��C�:�߽�Ǉ�uӮc�3Q��3������'�V_����������[���[[�:��3����}<���U�n�6�e���йѮ��	��d ��Y2�x��a������걅굔^��K���_�'�V�b�e��k��c��ǭ�#!�2�`��zDUR�@��v�����]u2�J����Jm�HS�_+R�7+��+����R=d+���"���F5�R����6�x͉��l�g�ª�����A�2�G�.>+!�v�=�fLH�T������e�j"|p}f���ղ����٥0�ݜ�	[�(�]�@�d�=6�3ST`�@�oUh���Ν/�0���J�'�a�6�	���^��G�5��/^�ɱ��e���� �G�����9�%��0Ѥme(��DDCC�o��l�䁒Zܼ�[�s%3��b���R��.�|�(6;	}��e��N�P1۝r�C'�,�+�l
��Пw>L��A���y��ܥ��~4`Ja�Ъ���������JE�8���d�`�f�H�м�L�!۳9w�$�~W���:lzD<��h�&�lk`��C�ސ?�Ώ���ͽ}w�|�/�Ag�*�E���W�Lx�=a7|�)�K������s����Չ�N�PD#�r`w����3|�N���Z�%�1��y=w���Q>��r�L��Z#��A��$�?q�q����I�����_H��˵��}룗Vź�Mqh��D�o�����wabu�bwt2Q_Y�,4���V_��^��z��S;�FhS���
��;���萷�5�� A+�%�EWS���i�c�%٨�KyS�t��p��֑M�K&����egR�ۯ�x{Ӓ�?��%�z��J�<�y+�B���5����a�!�CB����78���y[/��B�m���E�æv�	Ho�Yْ\�& f��r��g�ϥ&������T`�}������&H,����G���{��a0�~���k+6;T4�~�N� ���(������F�}~aN&IN�N��O|�-0^|�ǆ��K+���ӴP�qxL�ƣ�P��~K��u{��m��5i��I��/�6�v&o�҅aK�l~�]{��w���<L9n���<�%�ʳ<|:$Nh��BAf�_�A`���{7���9�C��T�u��`�>߉0첹V���א��y���2"�����P��6^/��I���]�a���_�5	��a]_��;�7�p�?��}W�<�V�aЈ}�������>�����,�=UEr7��\�:�(�J�ד����1.jNL��Y�Ճ��׍�&>����a�G��¦\�-������:ۍ.��S~]E�?�K4�D�h�S��:,�qz�tRܘԬ2�ڗ|��'̕�G6,Yc&�j�RG�?X2hI8������>9���<��#p1o��(�&��.�]i�j�%N�w�/�˖(�8x8�RSԕƵ ����Q^��u���d�A���^�k���}V"RS�8n����z~�M)�M����ď&[~�~ѧl��C�ȳG/�N�*�Bi�x�܊�9�D��[��ئd�g����S�5nz�/�z��8���<Sko���[�յ?{��WeD�2����(�CKt#b"̵���\"����J�d�&���Vg��l�j�3e�n��)��@�'��^m*�Ϳ��Af4�C�M�<?�T��F��?�cNf�O�ʕ:�;S���9�Ц�Ҫ[�̗6�.^�u��˃��� ���!�	���X��,/�6�+��6��ɓ�T,O,\r�ND�<؅+�{�x29or�ϥ�GQ���ܭ�h��M�oEU2�����?0�o:���(e�#��x;����rk��x��sxy�Ս��/l���⛲3�DϠ����29~P@MXQ�����xNՍIu�y�������G�k_��e{�|�����yD'��G�<g�W��a�Vl�AI��e�,��v���2�����H�V�)�q��I�&����Umӌc�7�5+(}��0����M��dYK}�n��ni�"�f��/��-�*�'
;������?_��������˘.���A�:�]�s*�\-����u8���b��v=/���ͫ���o��W�����0mB�P�*%����F���� ^	Y��,>�bdt��r�c��bT���|��i_�_S���ʋ^bD8�c���:p�Z�Rғ9�ወ���T��+խ�5�k�_�|)��Q�ns��9�Ƴ �{�wl����)���T�/d��O�ޭ/7���N �-NQ����ֆ���$��
���9[��?r$B>1*%ԕ���
1y��+ˬͮ񴿣{���s|T�S _���^z[���m1P�)���}�(�c�9=ͷM��jͨl+��h�E%��q�9#P7ROjE��кȼP�K�Sz�̜���pu��Ky�`s���@��8Y�R������HB�!Po0�m��?RK�9�m^<�r��ܛ1���>~�Z��{���qsi�y�.Y�ɪ��Z����������<�.��fb2��OZ3�&�KVMfb݅�k��-i��jrr��<�cf�<eI�I	pEZ���~�=�K3n�����*TM����d��1d� ��t�/���_&��?���_�{.�|?`���T��t�c�*�$v�;3�:�&�5�$�N�YL�\f!�������s�'�D:�Z)���ɻ=�Uv��J|Kg�+�{�`|�,�K)a���=��R� <�g�QY��M$�<��F�&^�e�"���њx닣����p�q�j��ޭ���Ⱥ���?�փ�8@=�o�����<��qj���F���b�J'~���/������?Gz��r�g�����~��;��/SI�m�7>�b����4��
q\�����Q#�v�u��{1o�9+�b����*~�7vU���4�+%ƛy� �i:,�6��ʹ����Ζ���t�p���>~%~�{�4f������"k~�������q��[�\*7[p�;��&�|�����|Z�Vӄ4�J/�Fş�ق[5�nl��{�ѱA^�_\|k�p����5l�����)�K/���e�����%U=a����jDK�X��a6��n���FE��ؐ��r�/kI4�x��E�ӥ��z�v�{\�݉�@���JY����Z��U��#�){^�bx���?Xם��]���`U 6���斳�t�y"yԳ8�_?��"[�;ɉA����h�_���F��)�㨷OD�D���F�i.�IO�3q��q����lR����������b��\�g�X~��e�H�Z�`[�DL���"p�ܗH�%(�bO�y���u%�͹�#�>��`u�n�f�^d�={dbaO@��<�o��Pc�f�oި����*$AH�,`�G׵n�J�ɭ�UPl�7߳�/{o^b|,�$�\^{� �C�%��{�6���R�1Omt ��;���f����&�WͲk�ӳuN�����ݍ��
�۾2�t##�����$�Y,U��N�QRڅ�%;O>]�j�I��J����4N��Qh�#vʴx��7��q���,$���kL�����̵l~�MM;d_++ oBUQ�Z�,�����v�?�6jy�9�~�*��gO.�N�8��r����N5�z[�v*@�''I�گ��͖}�!��M��^a�Bu��%����¤.�JC�N��������|=��T�+(��+fZ��,�)���u���F*4�Y�4n	���$m�O��݄xx�^[5ka0�@r��q�c�,Ɛڏ���^�*��'^�!s�f�X"�#:;Y.���h�m���i��T���Qe�+U֣R�:�������! r��XU5?��m������".ë�>XH]Nuy�$ޥ�w�մlFdv��&;��D]�&ɅTs�<�����PM�������܇rV��+R>L�g�N`��8�@T�3��g��[H��Y�F��� ��//�(7fu�ĵ�E�W�,�eBH!t�<�4��'gq�Mq<V�}XU}�P'�=�ţ�����xyX�!����W�}���f�5-x���ϿUhfaMx�Ⱥ�tU�/�&��`�Z�b�\_�$���G�������-��W�x�i�~7ae�m�l-B�kz����y6Z����}dH:����]����>�τ/'�b��5Z��\����������Z����J>֐-L�7g��M�u'�|�+��RJ7}�u*�jۓW�l��!��ҳԑ�+��CJQf�U�8��w�K�65M���� �:�&�tɻ����>$^&? �I���u�!�1uf^M�{�tV�b�\�Rn��8���' �Kȫ���Ug$��ֶ�|�TA�'��"o�!�\�g`����)N���������u�7�+����3�W.������Ao�ͽ�����t?`S_iu�&�pg��A�Bº{��w7W��?n�y�n!x=i�=#W�����<�u�YV�!NH)^Z3�0�׋�;�x(�6�+Ӻ��[o�Pz��=�>�Rk��K4/���n���=�	NbYsL=?N귄'�ʴ�6����2�imC(g�g�b/�
`�	q�K���Uys��J�űǥ�ٿ�H!7���9[������/����.��<�o�w�)"����x_.4F׽�?>�f��X]��{�������\\1+���-1�n_�IJ_,��}�ɫx6X����_���|I�>��uN�!AW�< f�#*K[t ��}�v�'q���U�S�8N{?A���-��_�s��#�T/Y����:��<N~&�G��w�ZI�X�Έ�QO�	&!Q����s"'����op	�
o`�1n}�YQP,?ڴzlҴ�+S��a��P�����3�ь��Me�=�l�����UI��:B�[�S���V7�[Sm���,��p�ϟ,;f��o�S�X��5,B`�~�$�Llc��A�vˍ��t��V��ȵĺh+��Y)̂� ��5��t=�I���^�U)
��U�VN���Q�=�f;��!�:Xx�q�G�λ�N��N�Ō���rl���UB���v�B�]yP)H�E���ȩ�D�'����7���v �!�j���m���PK��ME�)qy��1B>�hjoXGO8������t��X�KXxIU��lF��,E��iy�����wsT��9?�0����*�;�:ǨΠ�M&h��ⶼ�fƭ���X�}�^e^̽���͌���N�Y��jǷm��ڸi9����YHϬ=mkM(,msk:������n��ék[=7�(z�12��� ��[������y���ʤ��9$��<r�G�Ļ��WY�:>�.�y۲kj�F-�2W���L�~���k��� �^�����<�cC]�gFk��_��#M���7�����Z7F�i��YH�ޛ�s^�Sh�E��U��\=ǥs�0�8��
9.��-�(�oM�{MN�_�2twq{yT(#tlf�;�M\��b�B��\S"�w�s���\&����M���I�y)����-'�&J�{n֢��0����lxH�ia��+D��8Co2,���/��p+]3�D��H.~j�؍��2�t��"R�y������ɿ7Q��ܕu�nlF����R#�<g��w�[���XU��]
�r'ln�ɪ��v��������� w!,��;n�z�� ����%f���&��G����-�ö:�,82 �h������IѭT�O�N�ObF1���:Ŷ�����ϛ9T��`�\"�[��K:y��(�8�T�Ɉ)H%����i���O!��[w�&��nq!�̻MW_��8=	�f|��>�z��8�G��z�̹|||S{�7��u4�X�O��nP;�,�k@w�����G�҄��s����k4d�ac�1+�J�wǏ����].*7$��`��ӳ��L����-D,�+u$n�����\���u��[V4m�(h�u��\9n���C#w��un��Ó	j�I��_0v,�M@�.�-�C��@fU�Ӓ�{�{]����O��J���'�����������K� n����Y�8O}�p��V��:1����G� �=@�h޶�X��p������-�5u~�{�����(�]G�焨��HJ�P�f��R�s��`�_��t�K�Cv�)q~� _���8fs2f�x�)c]���J�d~i��Ѯ�⷟ds~f����g�	���]��-{8���f�m_�+fT��9@��K��{9����A��>m����^<97&]�M'�+�Y�K�X�]��R]�;I�mr �@W>Xo���Ts�ZT��l�6�2Cφ�M|�Y�$�*�;O�R�醎UT�~�Tv	5��J�?�ƞL�ڨ��{�Scl[b�׬3~r��
�_(����HMS�᝿�.q��mZZs�Ϊ�
��A�˧�;���Oʈ�n_4�nooB>��&�����9/�<���۶D�� �W	hq�����d�bfxU�&wmAM,�I��?ɥ��l�P����E u��-��ļ�h�KQ�y0��~d��s���T��̟-Y,;`J��"��xo�쬖��� �P�Y�9��Nέ��P'�Y�aO��U���������J��а�e�sV]N8ci4��L�zuj�7"}l��[�X��κ�W ]�d��V�ۼ�n�@&����ą���F���d5N��b�ܠ�l�,����ߩ��φ��Ϣ�;aVo���)^3��x���ӳ����!đں>4-ķ�a`��F�:��o�F&�Ǘ�ڠ�}���ɋ3\2��)�8>��x�!'���!��8�#�)�Ŝ�gѦ$�l��-��#8u�� ���O����
 \ ;p߽�4x8�ǯ��ӤUE�)��`��N�6�v�}L������z}���N�Ivhi��H�.
���^6j��7�*ǡn Ȕ���g�(��<;g�k���=+�l7?�s����@�h�55�
ǰ��C�L�uw��;/I6i����h�3�ltޙ��G�~q*�
+�(�M���i�ǃH�J%��r��gM@����Ɣ�~{�m�u�%Y�0�AV$K3�T6F����;�C�l���G��w�_���� {e���=N���ׄ4>��sͨ��07uځ�����OSk�7�r��o�{����fp�) 55s6�"��<��*J��K���
Js1͜k�q]� �ӗD�䌴�����n�c�g��� �#_/��̼$^�ڳ�F�2�C�������$�n�Q���>���v�ȼC#H��z���#Vv�k���6�_l�%�h	hx?7�`	�Tc�$����0�����|	����˕3�c���8)���Mz�kU���Փp/�=�-�F��3���Vs/���9U�)��IaW��w����N�[�Q�9�zي`�aT|�Z&	���cT��gL��ʻG��gA�
>]_X��k�)��z��ǉv�>�`B� >�=������r������#�"P���;3�����17���/Ta|�����iӪ��($���͇rv�����������#*HU���5` ]�d�,���,�
��.�S`_�fa1�gϜ�ʵ����{����f+ꧣZޔ/6�����K�����g�Vf�v��gC�{sr���� 6��_��T��1}q�O<��`�@��3}�SРki�h�����%S��5뵱;�O�����yCs���_eq��⎦$V�RNם�v�����g��$�_���~�׿��h3�cfZ(��/f�.��L6�o}����8<eDZL�(}���<�\@�N�o�OQ����-X˦�.4�"��.8C�s���(�ʅ���e⼝s3�x��~��p����va���6�2i�>I3�8�B��uG��	̃M�<��wث]�L��Up| 79��ϓ���Im��%q�����1�P@����@��t���K��F�E�%=���fx� �3c8:T��j�T�Ӻ��тq�M�K�����S`e�����S�ތw�/�i[��ރp~����&SմM�ͧi)_/�p����Mh��U�[p�]�d��^�U���D�Cb��S�Q �?~}�<�%~���1Fҩ;�kpc��$�Z͸�w �X�[�t\3����	(.�O�H�I���{�-�f�<��Щ��Y)��H_�IVc�ؓ7'��ܻ\5eLc`���8�櫮�xS4�I�ސ1��Sya���K�� ���r(�T��$�
hA�i�[��|��?'�>�:(�rId�Օɖ��}��g$[�z�>�?J�
�6�����2�C�H�CDt_pL��'8:d�FU ��cw�-�6��� ��" �� ��Ҙ���T~��4�\���O���<s`>�{x�Λm[�łJ���}!f�Io��7ȳ:T��2u�����}W�b���}-vMR������_���/�>��L���m�o��H�)K fY�����h��.S}Y��>Y:��r7#�}��������W6�oꏇ�Z�|ju7B��o.��y2k����(�xDp���؁I47�tݵ]��;+M�YBK{g�Z�ߟ�&�N ]�zׁ�	���,�03we�wߕ�t���'�+5M0��)���ة���v괪Nѥ���|6xr��e�Qy9�'�Z�Πԙ����6]��pc�a����n���?���]�y�ǅ��z��_ևBe���l!MV�Hѽ�4�bL��5�Ĥ�jL��h�xM��qe�oC�1o��ڑR^E��~�{안倳�ϟ!??��:I��=]ܠ���,8�u�9Bż)ć����J�#yEѬ<�q��G�j|�� E@�7")q��x-l5UDb�>P��n6Nb:(Zr��=�d�-��_!�=Hy��Ý ��g���.�O��ѺQ����߯Q�7Q���hh���0���$��fϵ1L�*���޻{}CY!�#�oTK���+���Zzrp��kh�JFL����FF�h�������=,}�F��B}[�I�|�i��bCB7�JŅ�&VdI;��3/r������(2��l&{�Qe=|��H�_�p(ܘ���Osû��K�UQ�H�o��|#b3ʹd}0!�Pe�3����Q��-��]��m�������1��}t}�D�H������?��H���1��b!��^��J�����Y͹�q��7c{�\���3��ͷG�N`�玵�}��d�j>��$f��)�-j�ri��3+R$}��E������Y���P��C~tj&<ֳ���N���~eG���]1�9�V�6��οv����n�s��>��)��hD�F�k}�A�A��%p�Ͱ�.�J��+9c�Zۣ���l�N��!��}eञ�S���J_��`�Y����1�Y�~�9D��e���7�]�8��}hĞC� ������Rk�g�?}=�:�c�z�b���Mb����k0��T���v�A:�5gS!'}�5��6�j�J�N��4������4N)�����n+�i�����}ZRl@Cעr�<؃mK��↻�a�M��3��:�T�n�~��JЧM9����r��Yg\���ˬàA��\�OS6sh�&�K:���A'b3qw���r���z���bG��%&�*�n�(��R�zǣ���mR��6J:��C,1x��S5w�34�n��r#Y�$k�M&oVԝ��p�+.R���Ԯ���Ɂ��s3=7�}"j�WV�n�3��M�O���Mȅ�����![勐QP�vщ2p��Cj�,K�g�A������<�jO�X�y��J0��j�i{�7�:�������t,��R�v��~����6"z/޹����S=~ĵ�Қ.����(�Tӿ��ba�j�����sz�Sl:;.��|��ـon�������vV��|&��Z����_+O|��K���1���u�4upp��ضHD��/�6nm۱ uL�3(��@I)�������<�d����=/��u4?4��l��Yf�0a�[ZЦ��e=0f�.���Cʿ��J�����0�.6����ؘl�A������<��	2y�0�n�>8����r\�Wc_�J���cO�_�_?�%R /U��kmb����I�:�/���{�!���Ū� �!���OY�p���o
"�_w����F��3�?���`��[{-X�U�9�c��X��ܱsif�?��EM��$9�×�&?���zԬ,|�N������j�UO�T�.�/5��ԟ���.N�_���5��q�]�F�&܄N�Om�k�An����s^R�_�o�f!�A�Gכ�-7�'(s�	Ƶtn$��܃%n��/5��E�Ԝ���D�Z7콽uWsa �R�ݥ�^�F]�t��§�-�ҹ+��K����d� �@V~~���g�H��M����o��aD��	7�R��R�rE�RZ�:z�}��$�>�lb�oo��.jW_����ێ'XKBC�߶���ǌ����X�#��KO�����*���(��`�W�"�?4Ѭ`DƜ"����,��C�r�˜jN��/���_��k/���Ӝ�m	�sߚVEy���G����x}���*�q'�яVZ���v�����JJ�_w�i��l��T�%��\[�b�q�k��T#+Ʒ�ʏ���6������g-7���Q�g��ݸ��ֶe��K�:��9Uuc�]G'+.D���.�d~�J�ʏ�i��+^�9�]&�|��C�q&��`L�	z�L%�r*X������Mo�qs(�l-��H�#�=���!ިF�7R�@s84߶W�K�2�@�񉃝�q�Y��v�63�y@i�����	3m�@}wܰ��7��/._��dՈ�Ϝ��btD<	c��Q��>��zX���5)?X�ճѫI�g xQ��:/�="��7������bۍ�Q��kȴۯ�k�������3v����c:w��6��P���vj�P�f�/J�[84�8��f\i,N,�W�Sx����j1t�*@Wɹ�ֲ��RI��?����z�ded�.s�=޵]4d�e-���U~>=?��k׭�����:P"К��L�j�@�G)���>���q�j�M�W`�#!�5��z&[�l���e=X���N��"Ĉ��M�����k]��#��A�[| RHO�;�f\d�[���߉�&J<:q�K+��hu�i���f��hB<�u�g�(�Iż>��|��@�`���_�崾�!����C�L���~�"���3��w���2�ԲG@]ܴ���BƠc狿D�u����M����d�g����Fc�t����Ź�ܳtv�_��۲�c~����cޱ9R�ϠĈdN^=_sb��_��e�m�z�آk6�c �Hm)�>J�s-�MަǼ4Yι�����Q�V27`�-I4��#��M�ϵ5T�^�N��N"p0�b��p�l�ztcUvqO�rH���Qa�|�u���I��VP�O�J:���!�ti���2敃Tam�^r��E	�L�1�~�x%�R������@�p�O��0�r�^<�A@(������RmV�����Ը}$ɜ�򾎱�O��U����)�v���}OVx��? Q��z��m�k���8����Ū���DN�/2�b����=q0�wZ�`}�����(�u����-	G߰�7Cwݓ�+��|�?L��M|P�B�a
/���(Nq����gp;����D��T�i���1a�{}L?$�L����˞k]�X9)+����Kn�'O��&�,c�н�%�;]�9n�xC��g(��9�$�C���@p������28����Cpww���u�wy���A�=�n�Vu]3=7E��7�8\�<���;o���y@[D�j����G�<�D��H�e�@/�Bm�����g������ ��m �1���t�/P���r_u�TwP,�H9� ���X��cb�C<(º�:_��3�TG^*�2��fa�4K,�|�����y�4�����eufg���򦐼���3�!s3��5�3CmY�Rspqyߥ`��#�~)���"��}��nR�n���v�	p���M��IOC�]����S$|���9a[�o�;)�Fo�վr��Tf|�]Z:(	��^��N��^J��N�"��+�N�r
SR��1���V2W���ŗ���SElq��@������z/�Õ�6,዇K��i��m��0?�6n�BY
��Í~՜�/vAajZ�X���	�	�\X�~�����d	�}\�W�ww@xB�w�+<�Gbg���/X�̘���?u�k0�M����?zV���E�8�QZ�J���nD�o-U�6�'$$�'�U��C�W������!H�᪄������J�q��dƛ"����o�P�����c�ٙ꼚�i�;Y�r��JVC�AG�R��������6ɴ/G�� Q���l`֥�eL/:T7=T���M-`e3�N���[Ni=��������w�v�6����啽��m�aڟ��/=��5nKFY~�����i�锉d���=� z��OO(�՟�o�����C]����+�[�nJ�Z���$�xm_�nފL��+%rن�΀���H����ef���=�X�Y��V���Iǵ�4�,�)��	nڢfI��乄`\>V�&�~["3ߤt��sœc�#��.i�V抝 h�7�±�ԑ����V)��ȩq}ݙ�[6�����+���c��0 �;�c�����kCMB�7Y�5-oe+��B}�"��r�&���=�{��A��0��*(��u���-+#�
)x��[�xnr���s����s�?p�ca}˪aA���ypB��+|%d��k�WUU�D�*�U����m}���?��9OH���v�Z�H��v2X�,������"K�!*2R�t�U�cz��wz�'
J�PM�����~��D|������w6��$<�'$fck��L=��fʭnV>�_�h����S�*y4�R6�"V���y� N`'�8�xX���l�1�T�J�~���:�r���8��,L-�='&@��Bmق�5�[����a�LǺ�G/CN��pn�$�'ԯCG���O�v��cu�A7��)y,U�===���/�> 40e�j���K�/s���%�\ �2��>\l��H���W�����,^ƿ���O-Ǉ�߽��v��(}6�`�z%�+f��2���[�Iw�ד�ƭSL��
�Fo�v8��qv[;��Y>{҈05�dx�Ɍ�m�e5�l{�T��]bT��ǟ-O�'YU��п�����)��qq=��J2�j�,���)���Y��+���q�O���
E��5�7�U;uA�ݢ�|wlOR��� >)(+ؾ���oO�-��,�mqӨ�Q��_����<��C��Am�`�IKDL������,�׎���oW}]��Ov�>M�$[O41H���=�@�$��Z�L�֕C�#4T����!�����	�������d�7�4�����}y�p?[�H"S4T��)$d�v�����-���-_��ߍ8˜��lޫ��n�N�ɽ{���CO4M<9  '�^ᧅ���VJ8�v��C归����a��M��Ɂ ?� I�����e�B3���5��*�^=�@�w����=��veT��ؔ���*U	En/íc��߭�������cJ1��[t�^��u�f��!:����U����W���kVW��q�cd+Z�1�.^QQƕ�B�HV>�O�'H�I&^���c��afz�3d�Ř�����ў�^Zff&�.v��)"�JQ�]��������)��q��9���X���獣��?����&BlI �DdIպ|���?�K?���]� ��u���g=�������_�����k���vʎ���_�C��QP��;P�^�|U֭k�A�>�JV�H�jG*�:��qJ�E���+al�F{�Cg}��#|?����.r��~K�)��cgɌ_�.v��]��f����l�eZ��T ���9S�>�(5[�L���)X�:�u>h�fK<�=�fs�Y/W�������p���,��!p8GN}Jm��א8��ZV^�׹ ��NסI�&f�˿_��|3���?dٻ-0�����H��-�Oӑ,Zҷ��ٛ��_R��`�[��;��1w�!'��*2��u�6b7�H��}�l����[#�����Ox	��v��S^;u$��S�A_�Vs�t<rrr�>��X��'~����%��Y��z���o���˩��S
�j����&=}��q<9�$���ϓ&���������@�ۘ�\䉇�*�J"Eo��e�߹Ƚ��{��u�0₴��?>�a��ȥ�F+"Y�A������٣)^7ѷ�r�AW�����w����
ߴ�
3'�
7�^Uܙ��#ٱf�?�|�n��,�M����A@2����|��=�ggʶ�ك�8SB�Dc!���
�R�{X�oZ���tGp5=�9��J��+��	��i��M2[�ښ[�%iԄ�IT ����7�rDS�n�T�T�3/�h8�˗?(�(���(�����A�pƽ�'�����h� [Tz�W�Rb^J;M�����%�~pe��ȵb���n��db�RZf����z�j]�F�DιT�.W��G��iE��=��W���	B�K̈́,�������d}?�run�����E����H��sA�ם䯚��)G�[����o��^����}���-t���[j�^����(c2���o����f����g��(K��F����g"�� c	Y	�η[^���Ě��^vf���k����������ӣ�Z	kO�/n��!�q��򝖌p�m2C��So�p���z*0����}&+V�+���2���YKe� h�镈wU�s5U�O+�p �Ge����¨Y�v�@�J��<!Nޢ �9^��4E�h��.���԰�zWU4Sw�qKc*�d�/����8l]$�!}�f�nc*��c��1��>�� �ǚ��x"�L��w<6>�@���vZ�vV���@�	�!�o$!v�Q���E�͟M�t����p}��l�ω�u�f��;��M@ajO;�t��� %d�ʐZ�լYF
02ڟ��������	��{|2x�w�����̌��ӗl9y�c��LX]5�R��*/-aR-��r%D�m3�>��=�$)#=������+X�Td�x�����?P�tq�ocZEW7�5�kLe^m��({����+��iM.�摂�Y�4��+�����Lb��*����W"��`F���r����	@s_ F�z������ Gba15�I�@�q\�oWNz$_�85��.��l҈K	V\��9"� q���'�!�Rk�k����N;4k��(N�
����wz�j�{g�ʂT؆u��H���ۜgA��Ϻ�����!���Iܱ�]�x�����^
f��^�z�tq���r��v�n��y�J��!cqb�e݁����t�r%�X��9%m)��܃?�L��%|L���xvNe�Fn�ש�: �N�����O�n�$�sD,�p�`�$�޺��ñf9Ɵ`��
�8k�z��f��{6ٿ
���~��;�H)�f��Y\���<�ԯ�5�륵���,��y�x��Y�+�R� ��N��ʌ�i0B-=~�j[�Pai�{��{s�;є�ĀDڑ�r�E�3E,�lz8�F���Sl�/Uc,\��I�ScC#2�қ�̆D?���q3��	�?�)�gG蜾�j�2��v�b���i����b
��?$=S��!o6��f!�[0�#	��%+/J V���,��!�c�&�\�!�o�ρh�&�#����-�p����Z\�_���U��f���!{��K��!���6Ƀm)z_�U�pUD֕F���X��bW��i)p�徊A�qπT��"�����w�#X�a�s?i��t�B��u�7Kk�����Jm_/����yAoCb�f����;��6�S6	��Um;cr:��쐳��oaO�␿5/q�;ػ���r7?���o��gA=[�Tr׍=B��VW�V�F�m�MM��
A2u�H$�n9�A�b��kAy/|tՓ,�/#���F��g���!N{���:��>l�X��?�ƾ_��׭���1�0�)W6/榭�9�"�m�_���]F��J)����DU��`K�b�����~J����ZQ�VC�o�ܐ�T��)�4�����3�'���qЂ?�N3�5X?���0���<dT{u����c��	<b�&:�YK��d����J�.���)����=���v��[X.�4�\aɴ.���� �@���EU��t�e)�,�EH4�N�9���6�޴��'�����@=��)�VT�t��%Fצf�=;�as�����˯o�N�}2J���Y�R�(�%H~Vpڕ��v����Χ���b�k~�*J��SQ;���y�.��+)�%E��P�[t.d����s�6���Ő`�%�2.�fМBV4����le�o�b>&������'���:1M�(�|)1N'��^�$D�s��B�WaI�f��ac:�8��q&9SR�O_�x�7�'CC��4���bGm	���q.���V����f|!ԹB�7ƹ�|��cT'L��+�ke���|�����I_Ȝy*���R-N�S���i!�i�Zt��N^��Z�D�����BI�96u�W�(�%w*��6%��m��/���̣�������6Ufu�
t��^�Ćt�[o�kG`�)!���R7��nթ��k������lߞd����(��/i7����4�Ï ]wYR�cO�!�!�L�.�-�l2A�t�[�� �k0�M��01Y|3��|E���!���Y����bQ�c��Yd�G��>�?�H�Bx4��'hRf��8��!F�X-=.3鰚��
�q\�;�-AP�_���U��T��J��L$�+��7=|�#4k�f0P�_9����G����Q_��tx���6�*����\�����1���WTH�Z�{yڼ��EϋL�$�Y((`k#cӰ)��܏����V���]�z��?ϡ�k�>H/f�"�Wc~[��*�)a���tKP�]���;j��o��x���(�
qt��+k�����}��<m`:�m,6�I�K&��:m�
)�b5�hd��:,f�6��A�a�K�e입;7�G*�G�ÍeR���j;9����:��8�9���x`�o�g�	�Ǯ�`����A�I�v��N��)7��k�%u���X���2�;E0��mͨ�����-�4ڦ��p��$����s�#���=�T4��e�X�;W[�|�@t���+G/�}a��i%0+=1o���V�m�v�V��`��gK6�)�k�=eT��8��b�A�w%�_�{���a�nu�+�3����"Gl(~U`YWC�Cs����!l;�埲K"��icp����-�M{QLv]�r^S�FI�w&������(l	�,���X��X
�L��Ri�F;H��`�6��s+����cV"ϲ�9k�i�1��>YH2�Hr�G�<0�Y)�J=gS�|g��Wl��xQ�7�XM��ၫ�Da˹��57�}90~/�oʎ-�?��T��Vp]հ�rr�^OX�h����b?�V����eX,H2�=�U���k���l�8�����M6��J	k�z���s�b�)�í�'07�f�IÉ��+���雒��Q:%�N��_\'M�#�-a~����b�UO�Y5��E�n5-� �y��U<��?K������eW������?��o��c�ˇ��^¢�Uξ9��$DdӇi%K�s�~^���5������S"��g���{�:��%H,�^��$3�Ήa,�op|�`���o��|aJd[(�g{[(P��n��>?��{J�G�\I��{d���h��Hn.+��l;c��wk����Qi������r۬�y�6�0{���M�I��� �aA��Ӻ
r���a�[�e�G��.�^��U���m���b����E��r��vp8�<�c��0�憶y�k��aZlK ɚ��;he�4?X ���|j@|��~q�m�4��8����v��V�y^��ƛ�����_�u_k��ǰ���+r���j������΍�R�3`>V��~��E��\6�N32uG�<��p }fou���+Y�>������ ;�_ɸH92 +7qC�'o?'ԭ���LCr���ϛ9z���*!x�tڜ�*kC�TF#�/M��1{�N�b����[R�N��z�7G��	Jcg?v�sp�[�޾��k� J+s���[��m��s�	-h�\
x������m.�I�n��ij����AJ��5�)�\U�����^U�>���8�E��lj&`s�Ҵ�.]QL�?��{
�L��`��+�C�G�$��vc�E.p�V��P��)��K_{��{����h\R�C�.�P��Su�.�_�լ�:��E��A���`=����t�1:�.hrcr�\ n��T�b�T�e+�����ߕ?�5a��3@�J�h5�&�@T�Tv?�l��H�SD�̓�_R�S�{�&l8ƙQM�ů\!��]G��1�$U���ٟ,�?�5Z1�f>���݉[�;K��m�uqz�����c��и�"�]���K�V%h�����'��V2�L��)�2��6��âfJ��f���,�n�˻�TK��Sl���w�>�bӊ���VU���V�R�����տ�Yrr'�r����p��b�|�33c�P5:�G9�b��}�����4Ht��cӔ [w����2}��O�$���P\{Ɩt~,��w��n�U�Ge��.��?�8�2��0j�j�����,>Ͳ{V����G���� �X�`Tr���l��f��2�1��v�bR�{��9�����,���ǋ<`wh'�F��Gٯ��pI2$�����b�\�l^���<��f`��y���fU`�-�k�;����s/�a�-~]2_�©$'V��t��z�,��#��:#�EU$�Ⴔ-�*ط���E�;u>˼{	+�x���(�٘�R�fF���7�<ǜ5�G�w��*\+hJ*�{d?5�|
ڬǬb�L��y��#�FU�R���m�w�[JNv������s�������8��+խ(�17�;�1p�f1��%�_��2~Of���������ߑ���ғ��[������\$d���F1W��qr�	x�����2go���v�*b��uӏ�Ί�&�'�ȠF�ow_�v�N�9,*l@M����s���;�67�wX"��
����p�!��ok�� �}�P�Zq���W�� ')�;xWF�_���ZP�ܑ��o�+�W$pBvk��U�̀@�l�Ν���Ч(����zm��jVĮ�k��N�T:B��1B5D�fo����h��'Z�K�_�M���t����rYIģ�h����*�d2������*i�g�a����~�vW��Om��a+j>t��Z}�U�?i���ȼq@G���4�)dk�u�����[���.����p�`��c��Q��\{xKl��=�ܝ���<78�C^)ZE����*�+z2�g���a���dܔ{R>��R
iFӎ?���܋%�J.��湲͸�L�3v,
��S��;`���0	A��|��p'�bT��#+�V�mߥ��cpW��v�Й�i�,��3�m6�͝��,����dU���#iTѴ���if�닃��?��u6�пBI
���V�<5'R_{ ��'��k����0��{�f��=�L>;'W��Ҋ��o�Z�o�q�Y"Oo��Pw���MP�(���ʓv��U�U-�'�Pg\ ��s� )1�ٙ���<]X�:MwE_�|����%?:�O��׃n'C�J�
|���j�qq,��sL6xt�w��ʛ�JÍ��}�t'��a�"�2�s�i*n�lq�`(�D?#��/�G��� ��>Z؟5svHkd�Z��n�t����T������WX!hbnqk&��&���)ɽy�����k5���)j���f�=;̇1���[V���h�/;G��M�r�!y�5k�:eGC<g�t�Mh43��
��_35�B����6�At+�z<��O�87�_%������v�B�X��v�q}7��χܙJ�9�q��EF:mS6bY�
��
���]�f���I{�f��[ �D�M��|�W��b� �-�_wT�.�Y�n��H/��9(H��=cW�O�UF�ҳ5wd����ۀD{a�8��q�J5��{ƅ��k�� c�5��դ��!���!��+�r>�[���ccu�!�V�-&ی���KS�'P�q筦�|���d:Ri��ا5���f�i�K5�ņ�	��Y��U�3�u�������t��c��e��I��?xV�lӟj0���S�VU�����/=<�O�`	�R��0�1(��R�����
�1h<��١z�]	�n���";#��%E̚F��L���O���������M˅Y5%����=X2���rmPG�W|���Eh���	P�N�Q����=+G�M&y{����NJmGKp5�T�J��G�t�	i!��F<ͿC����ъ+��
�I:��j'�x%�ml8���b1Џ$�h��s����4L��^�UjC^��琛�0=�Gj]��X;��ߊ�Nh�hh�E�\�H>@�_I֡o�W#{�1�F�ҽ5�?#76��h+�I���wO�]d�+�M�GQ�MRY���7۰��>�ow�|l���=�Th�q�55���ַ���b�S`�U�R?�j��^V|��)�.�S�s�>���
b��	����V���e8�<�埕gw����sNݱ���IpsIaqqq{���i�ɡ����ٍ�t_��IU�z�{�8�.�a[�2ywN��OƊ��o��&�q��TU���ĳ%���k����
���zZ0�aZ�W�R�@�4`PNov�V�c�]ߕ�&5��]��j���*�.�ƹ�2Wof�_Ʃ
PB��evx���Ʉ��s�)D���PJ��^�xȡ-<w��j$C9� �?O��+��fl��͊ڞ��>׮��7����tK��ۅ3�lM�Ҡ����=�J�vM	���a%��Ic���86��Y�
��)��J�Z��[�Q���Rm�����dN��G��w̠�3����?�T��̭Z��z��Çy�ѻ"mǦ��掘'��{�� C+@�v��^���������S���؟N��P�	���Dl�3�H3���8oEe�� �����_j��ާ�p���������ߔ��5�eѵ�������@�p�5D`�]�v�ݐ���u� s����5Q����n��@a̵�~�F����
7���X�jr�������}5���e�ǳ�<DҒ*~��e���в�������G&������5z?��L.�Y.�HA0�#Ʒ��^#�W������$y	�}��Z���,�F��I�Z.��ܫr9>��8��J�V"TiJ�`�c��Z����˽6��'�֙u�U�7�F���\�p=���Y��7J�9�C�ߑ��Tu+��	��^�=�I7��M��\��S���	�\5O���]2��ѩ���v���_|�4��뻤���w{b,:���q-OGM]� ��0�[�]���R�:ؑ(�0������%�۵�M�C�n����O��n�p������q�OO&az�Z<�L��!C7+��g��!�����TU,�J���[��$3�@�%K�o&:Z��ǔ��_&c*ho�^��2�aǄ�V!��ƒ� �/0����cp�F���^���:�=���6���f��03KFB�9S���R�r4�װzx
�ʬUjԎk��R�~���0�%��qL��Wo��n4b�$'@�,"
l_Y�}D�d�Y�A�ׂ�;N++�Y|I��lK^�m�>MMx� �����*��$_��"�Y�1��J�Y|ֳ���K/�Ȝ����s��;�m���I>��~�A��F�4^)`h��>[�h��g$��|���#�}�y���
�lJ�º�2���1F��/�ZC�rmM{�r��
w�d{#��oҟ� V��|@����$��6~))'C ��|O?P���E�"A��h��@�ΤR�b��D羴$:�K�о{IZ#���ƭ���b������WQZ`h�S��Xdi<�S�hoо
�;���o\�[4�mL'��/���;K	�j�w��� o���`�ft{@��){!��k�nO�U����dm��<?5�59��7c��D�)Eٸ�vj[���BD4>1.�����܀�v�nX�|�ꔤzt�F$�(	�6;.�>O���/��"~��q@xBQ�&@q�'��;m+��+�_���	24Ѩ=�r��	!3n|�6r꿊��[���DbO}�ԑ �5S���%� _�O�;v�|�N�J�&�|_[߀�g�5B� 3�3uX���~ ���T J��~��_>;����/by*����S$)S��M�aI���� Ěu�Ay7�H��Fm�x+�W���r�mk��r�z8-����Dsy���7��I4�#�f��F>�R�[�$k^�`W���BV��90���"˘����-[/����r֕wX��������F�-�c����(�z�l�����X_�F["���P���B�C;�y�"�"�a
:�M�g�p*��	��6�f:N����Bb����O&%���t0_�z�����c��wô�7q�����z0���6�Tӎ����+j G����	������7F"W��&�co��g��*�ێ����{J\u��:J�*��N{4�$NB�0�ȣɂx1���zK�/7��T.g����T����g�,������P������̯�C�r5�_�M����^ַ6��A�y�Ε�K�n&�U�hh���!�����x��Kt�*'UUz�P$><����S���/����"�b,�$�*h�����6���T�KL�j�HI�$ ���۝�H�w|+�y~�.J�W���hi�!��������a��/�2���e��o� y�8f�f�=�ja�y��~(o�V�h����x5.�9=S�<
o�h������%Ur��/Zx����^Nn&!Po|m0�eg}M�(m�D^ +R��REҏ�q^�� ,�W獋7�=�K��VP,��d �Qk�œ/jr���Ir8��D����Y�a�l�U�E�k��}~�8�S�5��t�{��^���,��Ӓ��QV�=f�>Q�Sթ����+���(3F��F9���\b^��H����-�X�Ɔ�����:�`�}�w� �eV6���p��5��ɠ�w�6iC�J�/��..2������pu�k^�=3����%Ȓ��~�g�>1�(8�� 8~�x�F��X[��_������'�[Z
��*0��|%�?���+�L��Ʌ�'	-l�^��8el�oTdXr�{�IW��Y�ژ�x�[�:*�첀Pw��&i��=����lT���-.�p��1.:i�G:� �(�Q�:e� �@---k|��cVC�V����hǵ)+���z�a��谰0Ef�W.�S1���WWr��0��ޘ6�7˭)����|e_�D�8��L�\������S�n��(ǐr��Z�r���X��6|���T;�����8�I�u#Ķk�?K������ߘ�y˙�� ��\ɕ�U|���"�\��q�P=_5u���Ѕ���B�������Nb�s㎰3���E�7X��G2����� n��;�SAOLP�
cc�{��"Q̆�&��:p���4iY�ƍ����a|�-��[�ۑg����^���,c~3�����uս	\!�\S�a;;_H;�j�""B�Vڔ�o[}L���:�.���v�#���Hl���/.�Sj ����G=��n��I8b��s.N�Ѹ�ovvv�~w�ARg6�J��%�K���w2@��p$��,XEQ�_��(F5|��6ej㢆w�����V�p	�0 r�x�m����]�/�S�9��./a#�%��Pn2��T�6g��`�CFA���@D��i����Q"=u�<<:mn��{�t"D]��^U�s9��E:[�#,�&��ҳ�����Uӛ#j�\�S���C�#�xp�=�����ߑ���A7]
�m3"��ڳ/�f�a��Eu|6��0�t��L���qd��ܝ4&��B.ط�=��^�KZu����*$���������o@AM�s��J�V��|#:�N��&��!e�c�.���6o�g������N����2�p�07�Ƹ�huS�hN�;�Dq�S��#��;�%	�@��2B�U���x�t�3�f=K�mQ.̱��&Noq��A����:"SЫ�k>���۽�l�s!8g���g���t�KRa�Ϡ�V���8�����s<Ǹ�} � �Lo)��'"r\��Q|�����7#��d����$���n�0J�4\��8�3-յw�{����[Յ˹4�|�QX�&Ȝ���\�&���t;�L1�I�{8ˋWJ��ʯ�ub�ݗ>7n�_��v��������������Hޜ4e�L|��:DL�m���Ŗ��s�R�誑�l�)�Dve��_��f�s��ذ9�e�Io���܎�1�.�z�d�B����B�\kf,7�i:.��6o��N�y.�[��2�RB����Uu��)���kF�H��0=��ӻ�N\����(�E�S�����;>Ǵ��N��=lK����_�m̩�CG]��ڨ�07s�9N�(�e^�����
#8�ؠR�;��ő��@����Y�
Ӆf��[�B�2�Ӷ���'�D��3�U��k0�t���WQ��g�M�gY>l����4}j���>���jjV!�3n)��W[7��bѳz��/�Nv�fsqHˇH�uM�'��y(VvE^Ԅ�����9�zt3<
�];����$]3�g_A�����������k�1����	y_�?5��1��;9V�%�IF�[_p6�E}�d�я�O���1�C2�4���a�0����d���?��Yc� �.�l W�jǕ(h+�0�H��n��\��}�x���ӹ���N�*֍6�&��(�T��a�����6������u�k/*���D1��Z�Iw��_�G��v=�x��97���M�S��q.|ϒyL�s�'�m	"����۝H��tW!(�u�!���R*+Iʟ��K�A�t�f��z�B#(u�/ N]��~!�"�z�[�<a�FG+�9)������JƆ��K>ξkM!L>Abܵ�6B�-��<��޽�{����a���X��oƹ��;)�I
Z�#҉����Q=I��N��e�˾�۹�t%⺠��d�-k��:�~�K����	��7d��'�}yl	
�p�����Gc�a���V$�Y��o�Iu<O� w��!]�;E�շ�j����0�盌fĿk�x���x���p����3�T����"��YL{�Y�$�߄Ne�Jx��.�/w�0KK媙&����i��5�ߜ����dd�'�p�2�!�ÿ���}QV��6�1���);����).X d�T�-9��	�&Ԃum�5�"��۵�^�o�B�MM�Sg,��WDY��KA�>7��/8��B��/� c�X^b<%���w�5W̧���0��l���|I[
���)��/��5zU�3���w�/n�T���Q\i��ǘ�����93���,]�4HW�s�L^���dL�&\��R�I���2�v�V�"o�[��\�ؿܳfc���Rs^v��t����B�1ˆ����d�!��D�#�9
���YH���gU�vu�Ky"�(Ơ�#�?���ő�Ʒw�_�;��N�`�@�]ȡ��Q'�)��[a�k��Zl�-��(opOc�A�����)ᔧ�7m�}�hL:S괰���=r�o��],�֏�xE/�-�S~O�"���~N��;���xr�  �k#O��/NCZT��S���.W�_(��(����I��H��e�����Z�;�?���_FX��Ǚi8����GBP���{�ь	hv�s�0�D\�hj��(m�x�L;D�.���%�$�rw�f�Q�7[jdlh��l��k��!���U��tC��Қ#i"�_�L���:�5�x��"Ke5�-�s7�϶��	��=o��m��_azn���#����t�5�Nc����򻿭������;U�0"�\��)��V�,	��:-O��s?�Hg��H��2�x�љ$��*oT~��1�_��iq��f���G�m��7�jG���}����-
O���A��@��:q��Z+A���_(gC��=IU��7�Q)���@(~�/��9�%�c)��\����ظ��B�kҾ�F�B��k%r%Q�!��Ł�������T>���B����4a����dm�V�Z�^_{�v[t��&Mb0������zGVaqG%�'F��'jn�H�����.9[�ZVt�.Y"n�I��Ϙ۱|�=��:�X�(������Av�LS�
�e�ݥ�f4!4��V�|}��a6�y�B�}%�o���_P��F�N�Y��H���:eh��5WM��?s�����~��} Y���7����*@�~H��he���@Ĥ�~���p~<�%�'a�O����,-�^\ú�V�,�R!;�4�{Έ?�B�dݢ>�9��KCx!�����8!<�;���:sׅ�*��"�kD�H���m����w�/����y��ϯk��a7��̻�5z������K���ߛ�;lك�g+�!u�#�7�>�g��_�c�ǀ߮]�)(�
z�f]�iLF6����Ӆ����Lӳv��*`��f��ʂmܿmE,�uݷo�p��ye�x%1B�>��}�Ȃ��� c����j���q`cC4���%�/G��F�A�����TUs�ʚ)EwuU<���s��R��F�Cp1�4�ȩ�2fw���"�7���R'5�f�Ȏ�.�y:�)��"��vT<��Wl�>�x��d����ӁiMl�ӹ��z����E�N�V,D��F`Bj���]�h��A?X�v.�/�Re�N3��vU�? ��Lv���;��^�����OK�U8��Sǋ^_eSa��@�t�RN��\�.c��m"/���1�H�E����߿,c����pN*Q� �%�̇���������� �Sk�k�����d,�����_�^?�g_��=���.�v���6B?I��E����9nw���8���D�~��#X�6��A5�O�������G+�X�)mh��I�X�s��f{Y�38�D3�b�A�����#��+1�v�����)(t�����wgEA짠!�'��{����� ����蚤7�>�7%r�g��_�|s��(�� !�K����_�o����`zx����X��=����}#[�6fM���ظ��an|�����=,�x8KC*T��j�&ކܾл?�q�7`����bH�;�od��;�'�����^��dr9��z� ��O���0O��.���}��'݃Y�2�u��<=x��IP����=���)e�%<z7�@��#����(o�7�tLP�Zն��n�<�������!�{4��<4��ֹs1e4�������8���K[~	5k͛���v���r�ѳ��)�u��Z�o�~.��^-��'������rt���tX	A4�!�ʜ��N9gZ�!�@��G|ϟs�~�y���Up,F�3�H*|�2���Ҙ����B~�H�ܮf������灿�yU&o=��p[��e_eA��EN�`k����f2��pq���n��^��)]�tS�*�E��;�2�k��J�K�Ӫ\�u��Q[�� Bl����e�,v$���A��cN�7܃�vh�Y��q���1]P��g_���o�7+�h�"A���������р��n��
5��4iJ8R��f�m܋U|��N�SY���-[�X¶��[L��7޴٤��*>���>�\��şT�w�0��G��? ~@����<�x�#�<޵���Ϫ�&�&�B�M�]�N��5$�&�y%�u������O 2��?$��.�̉�A�D���S�1|�=�!�c�EC�_3Q۳�wމ��,�M0��)\8�*�=�89�Օ�ևQ)�D��G��ȱc��~���$��ߝ&(���&�)'S��$���5Ƕ7J�&#�c��L4�jd�:#. ˲z�V���]�F�'<]����֡%k��������"7�*��-t�>vy�T@�w(�Z*��Xg�i�R�����\S���;�9�
��펂-�јp��@���t���l5��1�,�hh�[/տ���$e
��3i)˘[\��;��;o���~�AW�m��}x���pV>'��Ɩ�q�8t���MWפ&�� zQ�ޛ����<�Q��T
6��jO�-~q9ҧ������]f$I�����R����J��{��?	l�����H-�T�P�Gy��z�Z��'��g	<�ji��x�޷ٷ=7옍e,�ڞ�B-;7n9���>Q���֠�
��ߝ�M=	�F�~r�������U����޳��SPF�}���x��(��6'��C��vl��ի�X�_DabR{��z�1�>w�g���q�_٨ի�t�3�h_ޓ-�ܻ�P����ajJ�}e�[���$c��5x��mT]s�IP�uk��`e��D�]�u	LG��ʦ�i�
��j/X�*e�S���`�\�b�4�*{��)���g�ɭ�����b���vR[-���,TN@�q�xu>_���W�r� LLQC[N���)���-�+W�࣏����|/��>������S�!���F^�]wch�6�୸E=�X:��-Vn3O���l�%ɳ��3����㌾&<�Vھ�9ϲ�+m'�gk�$Y��Ա��t��>�މȶ��^�s�'��#�w2�o^�J�;�����qF�<��R���p�8>,w�p��ב�M�jD��*�<f�7�ɄӶ��Su��P��XK���0}سOMOЋ	�*a��0C�{���!�}�uTt��~�$����E0���K* �رS���޽���_^���Ғ��G�ڬ�Z1��(��τ|F��lؠ"�LlVO�!�� ��a�9���vZzvLȄ�Պڙ�E��|��	�T�k�>�Qo6�
�LFX2g_���cc��8[?55�ep&
��ppD��1l���{ݍq4����$4x�7n*L0T_��F�ra���4K���w��==Ͼ\�iI�>��G�i��ͷ��}�;سi
�&'q�'?��¢\���@�~��p��:����n���H�kb$��>�,
�I���S���M|Nf&c��l���W+_~�����;�� �:�H��2T������0���ȼ|�A�u�r�o�Ư������#�w2r@��]	�zv�m��ʝ~�����Q��z�L)ngBv]ۑ7252�A%f��<��^��Z��C¶l=a���K�>�O�@��غ� aO�b��mrc�=[�\ÝX]ڢ�UL�*x鯾��>�!�N�bu~o�{�H�!ya��?�0.���6�
ˍ3U7��t����M��1��L�9�5kY�ֱ�(����@!�6O����w�=�ag9�`�36:
�`,Y덺3{�l*�����OU���a.%�胾6Av�r��Ж�4q�h�ș8�:_��U�n��5Uسo��|a����7�Y~^Ė���;�9�Ɍ<��~xa�s�U�����/���P��~����x��gtOK����ߋ�;�.�sX�T��(��d�R����o�'�G����e\��]�!�9�,D���k<n;6:	.vI���={��j=����n�\N��.~�����/�����#�w*r@������i-�Q@�WA���+H>U+�*rC쭮�B�T��Z7,��@I�#u-�WnJr0�kc�έH[]D��pDrc_>�&��.��};x�u
U��@�v�$,�o:xG>� �����V�Ӿ8�����G�ɗ����I:x��Wq�{���c��O�".�:���_�Ҷ���������Y5�� =�g����8�2�J�xV%�:d衰����&?d�g.si�ꆵ��l$���ظ�eBP�8���;:~FF���+��M�;U�MA[O�_G~���uú�����]��c(�޾��v�F@�fe�a���0�7v�ʟXۗ��HҰ"����$�yM �ʅ�ĸ����>�s����ۼw�s�b����i^-b���z��D��׾�m4$���}9�2���'����@U���c�ڐ�j�nbs�V�2��l�T��J߲���IǏ��0�[��NF4�^z�p䀞�;[ww��g��~�S�eJ��*K�g�t&y��DǣX��B�3;�#� �-�̏��Tn։�Xޜ� uz��k�9W�}�F�L�P[^�;�b�rJ�k��#�b��)�[�'p�?���]���}����ť9�|�5ܾ�*��=�_�����ͿR�(|�C�7%C' �v�VA�f	{�C��U���v9
e��3�s�$�|���T�������{�^��:p�(̭�YJWVm�*�'8k�����ͭ�a5%�@>U�<�D��2�79т$|������X^�'��/VQ4	�26s�9���u�J��F������]�������5;�G���v�y�%\z�Ms�,��'���!��y~�\��I��
�V}��E���S��5(�1�P�X]^�E���*'��ʃe��9�=u�|ƋLi�Ϊ(�a��@mwB�W��H��'�~�lb����J�u����G�d䀞�;W���a����7�D���Z�r�,p��F�92�Ք��c-ES�D!U�n �0�y�q��� fUwm����#�{[���a�籶k��ޥ}n.i�z��Jr�c۶�<�~z���f7����_~������=x��I4dεC���Z<�a���g��~cCCf�!�@����9�RQ����kDbaV�M�'�:F���ی�1a!�A/��.װ��wa���W�6a�U��	�Y݂����[���~;��5�s�?Ε�d��oW1{�ı�$KI6s���2���Z��V*�	.�k��n �>~�[W݃c��j_�U��<��Jr��r���>�ݣ#�11��+�x��gГϑY��G�`ϡ��%a��vR��پE$F�QBo����%�Q�U�U9��V=�j�_Q�-�:��K�����y��B>.�qtÞ$?%IB��\�a����>P��ƶ7-����W���_�m�G�#�w"r@���� W�+C�*4��-�]�&;��P��T���f���9���I��d�v�FD��̓ Q�ʚ����y*�զ;�������:s�7�n;�{ĕ��=f�ക]���^�}�E�{�9���нzO}���o��YF^l���+�.4qǃ�>1�'>�Y�z�����/��=�����5���8G�������9��ҝ��J�5Y,�
ټ7�4�h-�Y��Յ4[���1�Ɍ~�EyLOA�����=U�F�8:�)��U�?�q�s���H�%��r't�	u<FΏs��\}.��41�_g��d��1I�3��q!
�6�L.a��j��ri�n߻_ް��|��3:RW�}�0��
�m,�jD0��k]���$�N��/����H�B+BW>�`T�+�e8�DnU��ɔ/����P�.	K{v^��H���X>[��#N3O~I|���*n�'��%�����,-&E�f�#�w(r@����O��z���D�Y[�u~~,�ˣ��	m4��M��R��$SCtT��Me�d����)��% �by�7[��T�;k��%U�_`:��{߃�����{h���nq����ʡ?�y��k�q�GOal|w|�q���w��C��³8�8��~�	�q�]��|����#Z+�(dFv,I�(Z��{܅��[�JE��
�QD0�.�I�j2C��d���C�T�E��ݩC�%	!��19o���I@��Ĺ��v�1�ge�q�0�@�1��:��u��u<N�$ ;j�ǶB����M�c��Z�#��Q�U%Ϝ��>?0Z�q�s��s�Lb������vmv�ٱ;'&q�ͷ1{骂�%����v~�<ym���,$)ȹ�.^�K��ߠ"`ި��e��QD��m(oA�*׵V�SA����_��ı��I0��:|����E���P����if��F���$&���<��n�0����:�XIJN�ʗ���+���g9����ُ��ª�砽0oE�/���n�X���gc�iS	N�%H%˲;b4��۝ �M��������ٵTbo�G�Q������my�+W���3߻���m� ̍�+�L4����y�!a�=��w�#
�e�'��kؾs��N<��Sb^;�
�� O|���Cc��4���o���D��?��.�ۡ}� ��j�rA@���%tF#3�
���<$ $#�YT�n��^A�>��/u��9���jo[�����u�8�ٺ�\ [��S5o�jw��{iq�,��"��Z,��a@�De:� Ǭ2�Ht���"�$+��v���n#ξl'p���{fJ�����͛qp�v,_��[/�&�sE��?tw<�D�"��|O+�/���d� ���X~�$&x����?��=�X�C�������z���u���=Ҁ��53�ڨ�]�|��E�^�}9���\�$���S����7���Pw�g�غd�+hut�ϋ��,���?Gy�,#�<ޑ�����,�c?�G����}��BMX�E;R�_J܈�Xn���+7~QDE�9˘d�Q����4J,Kb,7W����%،��u�~�^���p��~�qD���>�v,����
8�q�`��x�{����f,-.�;���������z�u������ڟ�)>�ħ�_�%�r���o|=a���������Js@�T@�T��R�l�-�����ʂ��y������Xwz��}���Ǚ��Q�s�~������l!
��.�={���&�%2�$��K��ju{6�F���|]���c�v���8
��	F��Ϧ�-�W�_ߦ;�0-	��{�Z|V�+r���l���:z�8��q�� g����G��4JC�hџ�\�WE�1�%�|�^}�~���5����Q-���@���5��X+Cc(�N�j+�cIP��i��T_���)����z�*	����i$�6��U%�{r݊�P؜��G���Dǆ��Q����v/��u\�c�PDy��#�<~�1�O�IL�]��r�hj��{�u��v�c��f��J�Y.�t�k���[�Т=:)�*V��
�.ʷ��8Cc2cef&��
�Y�����u�.t1��˨����C���Ӏ,���r��0���'��4�������(�����x�+_�Bo+�j& r��k�������x�����5<�䓺Vu]�yɥ�ʇ��$/��V�(S���<���H�b�g�b����2}�0��8��Ke�yPB�q�����`&�'O����d�sx��h���1ؖƒ?�����(��U���Y�k$Y��&�t2o7�w�[*�K����ju�]�x|��'�mt��\<y��${��MLm�Ï;n�]I�سg雉	��x��:�o��������[��_�.�jwEXyi���abcfnA��M��Pw\���pE~<_��|^���|�&���ߎ��%�s���*�ZA>=/V*I��5dW������]�N잒k���Z�k��?�<n��?Cy��"�<~�Q��ધ�ɓB�?؊��7+~QX��
Vt/#;,U�lq�[n��骛��讯�ǻU0�O�-��0%G _續ى:z�t���W���^&
e̞<�k���|]:��*���m�-�6.Fm�6�#��vi�j��N<�*�'q���jݫ�\؁�~�$^{�e|�׿�<�V��0=�u.4!#f�O���QH��hU�ZCU��+WޗNqm2X��9�z�'��K�I�;���l�� ��ly�	����>ؽ>X_:X�bl0�s2xy�ِVDd��bW�ą: ��	��rG�x*��Q�(����}� ���1� q�1�aM�Lx�XV}�����:�/_��ū��lq�w��=��Ks� �h"R.��ZzZ��5���_������/|[�w'fz����( �Q�0j�(�DC���v�1���zk���p��)��_�c���NC�Tj>��$�z�~�����EI�������w��;Z���G�C��zܜW.#�<~��z?Ә��Of*iYb�Q��?W)��U���Ҭ!I��GԐl��F+da��H�̈[�|[���X���T	wg���TU%e���*�)�Bd�f0E>
�M�<���Ci�^t��x��/`fUmJ�ܷG>����/��f>5T��_��=?��'��o}/Mc��8q����>�?���K˫r�m�v�����rs���{V˞ ��z�,�RŨ$6K�5,������pg��"Ǫ�q[*,�U�ƒv ���9����يTI؏41ұ5Ή���o���ST;W[+#c�F��wQK�췫ɹ�6����:U�i������y8�X��b6Ѓ��HW6W���al��v���
V�]D�+�W���Çq�GAatHr�e|]�*��[��Z�U���}o����0��/��,�}�n��K��c;1F��c���0�u
�!sM�21m`|j#3�8���H��$ ]\鴰w�D�߀��x���\����&be�7I|6�~���/ؑ�Vb�I��A]��'>�����<��YD�y�L�%f._��v�!�v�C;FʅBH��/�ʎz�ad�N.]am�9���;)�ݶ��O�k����zw�H�����jԒ���K��2n���%o�w���8�'_ö_�"*���)]yn�T����E�\f2���E����?�oHp��|���_������B�$�[((��/��_�w�Gv������z�)��n	��.�%����eT0݂�cf�K��:��"VVV�J�;�J��]5�	Ty^����(���'���z��ɢi%k�Fͮ�I�I"�Ԍ˙x\u6�Y� ی�(|�(P��5-;��2����Vb�P�0�F�,����^>��$1}��%a�%.��׫�cw��&w���Xx����ٰ��]�����C�� ��S*��Ԇ<���-����SO���&6O���_�y��\ŵβ��8l��w+l�nގ#���I�a8���c���=���0��a�Νx��?���Z�(m��س�s�Z}x�n{��Ă�[� �]��Z�?�?X����Diڊ��H�D��r1w���g9���3�s}\E�\+˭3I�h���LV����x�{s��(��
2��ׁ�mc��bQG�茦F��;�UE��;�Sc��9���&���L-e�x&%9�;skϿ���8J##rs�CW�m����FeX@��ß��0�e<���Q;������JG� ��s���s�n���kh^�Ŧ����>t3W�%a	P��Zn�	�hȇ|�]�YP�q���\Cr��ڝ>ֻ=,���{�h���ח��&���HS�ʣ�=��H�;Q�(�zfz�=s��>�����/sf���9�3�^�Ԛ֨[ٔ(R� H��M�����cｿȪ"D��Ğ�ݼT	���Ȉ_~����.�g�.�	�l
To7��q������uS� ���{=�ȉJu����]���"/..dP$T�U����z�Y��9�"EiAV��T�ˎ}��s�@�U�,[��p�b3ƺj����eD�˸��I���	�]�O�տAu�v,y�]�R�D�ڑ�:����38����\�ǟ����2�7/��� m@Q­����)ku��+�G��RHɢ=�����Ŝ����Н�L�`�ق=TF7g!1��P���Iq2ą�۩��u{�k3��wG��E#J^Kt-�5�(�}{�;�����sl`_� }`�lV�|,Eq;V�EQ�8������9:�,�R�L�ow�(K��%6��l̦��' 	yn7爹xN�W���l�h�3{��������D�6H+��b�W��5�u�� W�(�Ĥ":o�'�:���CWǞ?
m+�?�	*)�[��x�R[�ސ��m���'q��Q��2��QԆ�h��[�a�s��:���z.�
+��	3��RQ�������'z�]�R�I�I���K�����2@7EHV)����G�I��.}��D-b��L���8�)
%U�*d����c��'G�)7���:3r�K~�+�9�O��K�Y(�=)�[�~1d�XW�b,7���,_���ŋ���]l��F����m;���⭂|_/3}�H����ֱ�8��[X7>��[�p墄�Y���a��<�V�z�&E�q�UJ�^�xh�)bFZ6�������8��k�y�����ܧg-2T[�!��{�<w_h(�Gs%1��a�%��������ZnP�>� ���Yl�'%Σ,�$��4�5��=��-���v�}*BJl3O`�`��$�7獖vKnu�q�>���-�+��l���.aI����e-��F�����y��N����rP��^�aQ�Prڞ"��<��59�=O?�9���~�<���	=�(�`��|l_7���1=s�:������OсBxtMy����QT���YP��8��k�E�On#����1y�V��&��:1|#��zFRl���a`jjR��lݱԐv��lJ�k��9Oeg�5�Jzַ���Q�4�t8�X3��r�2xs-��9�G*�/�y�&: ��H[YJ�[JޜENP��1b�[*��Ї�[n�1�D�hx]���<����ƛnA���F�:x�;��ؤ���.N��_�yb���&�����<\�R�Iש+���qTgF��u��Q#S?/k�K$e�!�E[����� l�dVz(2	����{���cF2��"�K��r
�l��䨡=G�j�h)?�<�����Ɩ��3l`_� }`_��~����Hp���8~ʈ��N[��c�M�Y�^�A�w�'<bYu]
��X)��dӳ�'�0�ߥY�=��K�5�qkF�#�i-#��a�cOL�������C{z~��&'�ܰݸ���G2ߚC�V��%b�q}�/�+��!��uڨ�1��1\^����K�YH v����HL�CGp�؇�MN�t,��r��W�i���RE��&��`�5�;�Yi-U�k|�Z�#ASY�-���$��}i�	�=b�<\��&�?;@|,ľC��z�)s(�@V��E�M�TJ�x��zs1GSz=_f�G��΅y�LhF6�6S�c��p+����2��V'gd���Wj����'����G!���y��݅����q���*����H���#�vJ.���4�����~����+ht[� r�,lHo�wy�M�LpW@AuF@��Zn��{j�Ο='�!]?��V��.W�'J�.�VT#�����p�=9���m��I;�?����h��as��r`��m ��ڭfÔ���C���D�-���c�B�fvdA���3��6Bq����tS���5�R]-��\�n�+}ג��q(���1f��f�a&+[P�b:1��2�Μ��g���a��
}�BQ9c��0�b��11�����!����_���d�ȑ�l޽Ub���P�r�{�N��4}��:^L�>ƥ�WИ�E���e��&����䧹H���� ���	����u�U��C܎#-d<;��Vz�5=k/S�z�j�����<{]֏Y��	��s�T��H[t�_��xMجD�=jN�!S�L��eG�st?�K�~(_$0���u�,�P%pޱe._����"����w�����0EI�g����KR�t�G�_C�m������Wؕ��Jy��.��a���r_s�˅�KW/bxr�[�g�7���߈���p����r��x�2�%&vݜ��N	�� ]:�l"�J���.=2�|^�0U*�.F��П!@5�����x^���|���}�6 �}����z��Ga�iq<�ɷm��R$tq�h�P�c�ŢTo3��y,s�9�}YN�A�{Ը�AL8$$�s�q�r�i��&��1���0�D�Дs��<�T7S�U�#��\F��a��øD�v�`m�$FH��&esf���@p`�����pk%��¿:�z�,-b^���k�n\n6�0l�V�K�\�E��������Y\�,!��ah��R��<W�K��.��!y-�$���lŪ�s�֬Z�CJZ..d�7��P����Z!Sr�UQ���63G��.yy�JqA@�3�����Tz�!�Z�Z�T9WHUovL�Iz=�`/`�p�C%�h��EL^�z���0�v�����0�q3Si"�-���!�u.����-pQC�8��_����~�v�O� ���~y/v�%@�;5"6^^����iT���qjT,��,cy�<]����c���k���Ioq�xpkc*."x���&X��K��6��w�>�z��m��Ӧ���#\��$����Í�<������k����&F�z9Z���������G�6�\�@G�hco���&m!n��(�A�ɡI7��r*CD�D�,�N�]\�m͹��\�(���nހ}#���I��ӹ�pP�y�VK��#&�~
��I�P6l-1	O8'l�u	����>�bG�+���t�<F�q����}]B��]�av����s����/�yy��*&����%̳��rE7�R>O��R���\�!�r,�*#fcv�|���~��������O� �JO��ihk�r��s��/��0{�J�C���;�N�R=S�S�M>�#2J��M{��\&�er�����l��P˻h�^ŕ�����e�u���#���O�%�I͑�"K$r��ډ�0����g������ob�� �Q��\E���!Z��F(�Mt�S1��s���Qo-�&�I�]���fc	�O���F�%�\<�:�/ۦ���B�g���v;>��y�������M���\L`�BvF��Q��/�=�|���9zn�-�K�l���l�4�k�3>"��m�k�Ɏ��>�Q7�X�S_�s�m��s�FV�L�c	 �����!_�(�5�XO���Yi̦�VXwfji��]c+�]�^'
Q�2�?��3�JY�1�8��6�/��%:�����^�xj�}�\��9a3x�m�n	�~�~n���W\��8��C��[8s�NM_�]*`b�F�	D�*�3o.�E����8��a4��� �eK_��_1����gr�W��U������L~U�j`
��c-�D`e��͌�U�⌕��".��U�[$Z��h�s�z�NM6�]S5vY�`"r����-u>)϶O�����[Do~���IMy�k��jx���î�n�>�J�:e�]�VR�<o����;n���yo��A��vJ0	d�ѰPrq��O0s~FFq��q�~�	Y1L''�3)���nb��H?�?k�k��o�C��/�#s-��3n9`~��J�����\$�u��vk���] ��G�Q"���R/��o!��G�ѳ9�4�=�y�?�0nx�����T ���6�e9��'1��[axo]3
9+�
���<+�^�Cu>CV� uы;2�����e�rK�J�Ԫ��x�J�t���%]>��ֲ�:�)��jY���@3!&�,��1�/c���_<�v���=}bRT�D��'���:3�V�6���'P���ſ��1s⸀D�P�Z��|�?Dy|����04?�ob�� ��֭��*�UG��@��D����Q��u1��JwS~���L�^��}k´�%�M_�k/R����>���b�~��ǃXtM��J$���8��2�-� ���O�^Ppr>L����b�qX�a��3g����,:,L�v�u���w��=��#�R�'��ł�PM��D�΁#)�^����������ŭ�<:���G�����v�I$�,ڮ5JR�O�'�6R�y�^Gj/\�>{���I�|�DN	1�*y*&�}c�Zg.�ڣu��\�(�����Er��9+��:��W�C��ֻƺ���Y��e?|pܴ^�U�%'RzA�<�ʀ��k���4����>����u8Ԟ����S��N�v�놦ž4�����""�B<Qo��\����n�n�f'!`��(TU�8<H$Ӏϐ��)Se�+�νI�����*�X��t%
bH�c�v��Ӥs�a� �ꋯ����������#�>�nW�����[�f7�_�o�q��_��_>��� F�^�KW�h.�>�;�Mb�����%ֽ�elj���:�>1Mրo�m4X���Vyb�9r|�j[�s�u�.t�
36.[*5��`�"�$[c�Y�r���")�� ��W����Lb�6��C���T9�X~�2��O:]��dʕ:�CE	쏾�������
� ��������"������wP,W�+����T�?}�y���_���6�YED�-}~���R���!:�o����c��m���(V��9kn�t�u�O���[��.�Ŝ�)"v*X;��������"zgQ�&p:�&FrC����*'@И��f��r���q�<�xT@���M秇���V/�����hir����<�&?�x��d@��b5b��s���v�$��{�=�U�l'��h�򈑰;���<�XU��$6�J��:�HE���6=�4k��Q�+!fd�r!�ښ���!-f���L�k�j�� ��\$�Je!�hydZ�c�70O�P��0w�r�Ԋ#)'0�	��"� ���Wp۟���k��ۿ����EJ�%��ѱ�N��?��{c�֡J�Pu�������,�sO`[�����8��hJʡ� �S�<_���2a�"��Cn[�E�7��ٰ���:W���3�J�"��%/�UѳĭX���P���H�U��>98U�"�d��CN�q"'�37���Mb�t ��߾�>�8n~�!�a��y�J��CR/9�p�r��J��Eo�>�"^�?��W�^w0L 9M��%��{�(��y6����?��.\��������Gh��������0����c��s�G�1��J �k�?�NAg�R����9!�?.R,��-I�,Y�,�p\�c)��x�3� �{K.���M�sva��X�e$�y�����別�{�lz�9l`� }`��{��9m�n� o2�	�'���p��
����)Z� ���h���h��*j@�Q$-X]��@��f&�)�wh�k��J���q�D���M��8G�!Jh�簴I/��9�&��x�0.0L>����#rtx<�ǉB	������!j;v����p���p�׿�����lH���
�O���wi|�S1U,�K,x������a��~Vd��Z�|�1n�4�U�͹QH�D%MD^�LMӳ��;i��_Tr5lGK��ϸ睅elS���B����:S�d��6;!.��r���'f�h�o6�Z�|z���x�������1�g/Rr �D�Ҁ�=qd�l� yl���ՅN�=��kx�?���lԉ��}[��j�U�������=�Ϝ���CX\�Ǚ��*��:��w�8ĉ��?�%-�QZ$x-r@ɡ��q�,51}�<��G�e�t�Ds�K�74�Ob���5IQ���''�A�_(a�-��z�~	��7?�����6��!O�>��]#��%]�mm���t�J��V<�?�O���d��v/�eN��&N����������i�;2Ɋ+�5�5�'f�cR#�fW�/�KA�oyӕi_���-�ҳ��`���M� Q���9��jͻ.�א��JHĐ��G�wa$��RSG�x�t�1F7�0�[�{�0�&]�}{	�tP�W��닳PD�G�1樋ݏ=�҆���ŗp���ѽ8�:��z�FD����s����c(_��P�J%LN��3K������иc�C΃��z]�ѥ�b�y[&�u�=�~*���O#q8^�r�"]"*	]���ڙ��q;Z���0�K�s� al����/`�RE��)��5l��` ����a�Z�\~��S��Ia������~Cr̶H���a�V[K��G��9�z���0��R,��s�͸���v�u��u�����3�Ås���(�"��5tO��<9���S0j%)(�sy�11u����q��b�b�3����:>��'�	ng1��B�i�&��:��]$��.��4}��ߌ���~ǝ0��t�t��".����ߑ�Rt`7|�k�q��(Y�}�f�z�v k�_|�aL���'� ��'��#���6m�qkf�lj���Fl�#�M%�M�u=	�FZ��}���L�K���Hz���0�1f�����\����א���\������
�W`�t�C�z��`��r��jYDR8j@�ѿ֜��y"XL�l�#���;
��,:���Z#�\@D����'�I�>�,V���ƶ�Ɓ����
��+Πf���������byns��Vº��'&lЁx�I�{�cM�K''i��F���.�
���W�2OocFK��Ft1��f���h\�NlU%����fJ�RI���'Ց�a��*���"Zn�4m��Ў�C?@�'�0�:p����?p=�j,;��{��:�~�g�yK�;�L`b����O�z�B=W��'0O̄�{mܺm#ʷ�OL��g^����A-�`�M���;o �kb�K	N\�ҩ���6QFjЫ�l�b]SB��-w,4�3pZ>&im�%���˨tC�t[RB��5:b�.��>�V������%����#�ޡ�ؾk�wݎ��9̿�܀�!�P��k��n�4�੒��@kq1!ǂ��墉S>�m���c@؟d��|��%C^=�ѵ�'�O�mUM΅F�>RD`�,NF�8&�*�L�9�ȄPdN:�̞MaFF֚�^�+��8��jUs�u��CNU_°���c5&����{�X��L,�}�CbumL�5a�q+�c�⌰�**�tt4/�P;"�op�FF19>����p�����O~�+��CJN@D�W#`��qJ�ł�F����Sm��U���@�ǆ�l.^��U*�	������v�Ȑ�H�HU�.�n���ֳ�pE����	�U��͕���E(�^,�õ ��E�ܩ��st�\���j5��{ny�Al޿_�7L,�0-]���qa$O����b�Nǡ�c�.��6^�����2�
1��̭�b�7oG~|/��&^�ݫ��fl<pvoކ��1Q��3`����/���3�����Kh����Ej�gd�=;&�-��/�y���#'(gj(�=9J�4q�Z�'��$���R��<���౱s�x���x�"�R#����eJ�������292,:h��օ�:�R�6G��S��� ��Tn��=ؒ������m=* �)qӈ�}s��P1_,�.����͛��Є)�ZJ�]UN�i�)B-P��Yn\�ޤ�ݔB.���R��������8��s�ݐ
0~g�0��H�SAp�a٘��\mϮ@KT�F|��i��	��]@��E�����HJyz(�vҧM�ji���H9��z�b	��ށoM��̇��˯��G��:��^E�D>@*U��r3�ʚ���?�hC���D@Z&`���sc��0r���-�6u��I�#���	�I/���hV�}޴�q�K�иaY���E4[���#%+au���+' +S��t��|��z�M�&Fe��GN��Ksp���O���q�Qr����;u
Ǟ�>����e�z[&����1�u+r�v�������g_��?��#�ܶ	 P��c��Wq��!$�����Ya����!j�2���Y��5:������q]Ou�~�k
9��^m�?y��mCr�W�����0W��qx�	lش	Q��d��m[:��RӗA8�j*��������C����7a��'�܃�c��/``��6 ����j��L#G�V�8~D׌��,�|k��e.�Y禚�EL����"�b��~�� _@��e���e[uUgf�*��_�\�� �Zא1�F+Ea\�-R#g&J_v6<�y�w$�~3��I0J�tZ�E,��<��`챇P��6�X`̓�rt�D�-v�X<����;���-�Օ6�@ibƮ�{�^@��\x�N_���it}��:�y�ǵ���(9��}��fX1Z�K��)n��A���s"�J4b��MN�����1zK��� �V@׾���r��$��:_Dl��v��m����زgJ���ػ;o�6}�vc��'ZZ%0Ը6�J��3�M:w͗@~���q��s��'�1V0�}&���0y�M����w���o^���8����'�a�$zAG~�,���oQn5��VC��D�ݖ^v.[C9�c�.��ˬ�n�B��X���]��͠˵t��:�\�s,L�;g�N�X�����ի8�����[߆]ǥg�y�0�s�<�(��������h(�KR�W��f��nҢ�qCO��ǰ���'��66�?��>�?ʖzL��R,�\y��O��|%���p�`q��p]DK�5Qmӥ:M�!q5�-��C��1�TO!{=����-���n��́`��s��:y�TDHX�N�4dؓ#a�R�I���љ>:���C�l�~�-H�F�d0]�JtvL87�c7S.�s�=��Ԥ�֜[1E,W��:� `���c�;�f�^��3�piay�J/B��y�.�{�t}���v�a!�,�@�Ȝ��'Pwt��͒��x�	O����w˄C��1:A&�Z ,��U�<��z�o��SS�ڳ�n���2R��Bq� ��t�p�X�O�TW��2Ն�$+�ȍF�C��Y\���`��al�lZ�2��÷�)��ǅ��B�%�Kk^����y�u�޼Q�����A7��Z@�b=�O�̈Y=�摼Y����i�����y��/���h]|Z�b��r
:mz�����9�I�E�G�S�7���p�����Gx��i�]�c[FQ۷�w�����Sa�9�����:nm��=^���%��F��q�[�h�� �/b`�*6 ��Q���){���IRN��~M7�����z�>��t�U&6��w���.M��`��'���B��� v��/�7_k�0�T���X��|K����7�ƕ֚�i�!9m8	b"��J�� s/�c�0e��z��i�gh|x#�B��=�jU飏��q �!�~J`�S���ˮ���j	糉	����*&n;HL�����D�~f�������_��*��$��o[��KV��<�vY�+W��qK+�q^�����+�Ιd�:��K�m����":����ҷ�ajvm݊�MSp�n�Ⱦ=p��T�E��2@&��팜1��F@�it�c�L�Ƃ[#i������ko��o^�5����:�RMb����]G��,Ξ�&Ŷ;�A���c?�Z�_��߰����a>�	��źRA�?�h5��D*8�/OT������2m��sxn{�N9�x�Z�l6z-�̲t[�,{�S\c���W�ֵM�Ņ�?��m3�ܰS�m��l �p�/�$G@C�>��y��9��?y�b#z�����Z*R���W���+[���d:W�[��xԃW4�_oҌ����I��g.��
8<�� еi�C�T��� ��s.t�u9?�*޹/Y�NV��)��/b�Z&+&ر෦�91Sb�� K�L���&�a�D"�^��jrb�<�%@(U��Z#N$�`Gj���7���Gp��3�ߴ��ڱI�tx:�W��b����q�����L39�)iU���r9���6�j\��Ko���b��eo�D�M���"�e�ȾWs�z䡢+��=?����G��e N� 1�we�"N�N���{��� b֝s1�~
��^wtD��y��L��H	c�tX�^C�I��CD��&��E�A�vȽ���2�xo?�"���p�y�ql��ĝe�?|�+�л�P{� �J�zTF��K��_Źًزa%rF��C��)��Q��]&3g�@1�V��L���%j�{�ɳd����?SSj���˱,zgfV�@י��sc�^ա{��L7Q[7��q?�]ۤ�3��#,��9�:�
�]��m��m����ۨ�82d�'��G�&ݰ��=��\gZ8�{��w/a`��6 �}%;w߃ M.vcv��SI�o��X��d͡rb7p`�-�W�����kPpΝ�������w�]t=O���V^��X�S_�+��B��$V�d~���5銨���n+�X�K%�ҡ��K3t=$,� ]�q������3�U�^�T�}�Es.���`�N�+G _�M{���	�z'N�r�po= ��[�+ҥ*�cun���lVuK���>@�c�P���9:�C��bl�v������(L#>q�^}=�]7@}�6|��X�p�B}l6�_�ȡ���<`���a�O9�����wa�߅F�ȓ�P)���R�s��N��XPVp�Q�Kt�H�
[jH���}sq����8��W0��i��e��^����wm�"4�@v��P�z�������^Ŏo�}�Akao?��N��M�}�6oG��'x��������9,�`Kn.���l#�g��J�@*B��a�MS�nҚ��	H�c�/���IL\(����Ӑ¥/~��D��-9�K���<��y`:��>��ˇ0w�$J��a��{���I4�|w���ψ�n����{��%��Z��q�B���G��u������� ����n�R��V���mD���h}�(U����6%�eTMb?Ej��VCZ�8���y���}f�����ھƖ~Q�\��@�ƅ
��ld�g(�7��e<i��`s�����e�ՙ�%%�&�2jU��R8�m�Z�/9yb�F���͸�zh?�%bӝ�>Dn�n8n@ᆽH
�z,�(��!K��ax���@ވ���z,玸',�C�F�X#ˏ��!6Yغ	ޕK��ߋuO<����x�o�n��'�\��2}t
��Vp��6a��#�q�ЇXC���6�u;�[7�p����{*'�~N_�=�(L$ܗιjN�p�Ŋ�I;��cXx���N!�8���:�#z�1`|�8��S���<���o��w��ǯ���-�(�و���۞�;�zᅈN���-4������֦���{1z����9
�$�*C�tR#�?M9�Z�:w}qT��|p�G�n$��0�P*�퀝,]�6I�DӢ㙁�Z�2���?Kk<L��4�F��ݱx���uo>
���T
*}D�|)6͋�}�5�H��oٯ���t��9آ��m��K�̃����ysb��Ǜ[I��QӬ��4�X��R��Up^ :��f@��۩_mb���jšP��'�L�tC�X5�\u�Q�B��x�bi�b,1j�#P�D �#X�c�Ce�>�����č8�+ó���C��i_��:�%�ޏ�K�9?,W�h2j����g�9w��A��;P�~,˴8�j�?�=��d'����p��y�/Xܤ�xf���b3F�W/��t�D:�[�<�#��BKl��S+��]Z�̑�8�.�E:~��-���Sp���2�36��ݻ1������h�������8��MףF���"���<tEJ"����<�\��(�؊���y��摜>�������)�W�.�D��uh	=�����{����K�ھO?g�������~��ﾏ�Sc�\L<|/r��tO���_<����߫������$�b�+2�P���H�B���30�s�^g��#V$���BW�^n��R�2 s�"�p$Ĳ�v�J�[��9.��;�H�:�n�����P��~�i4�Xf�\i���^R<,�K�[�~�~ی��I�-F��z�M|tם������l ������Z�	���4M���[t�(��$3��^��X�U(!O�5"��w[�{f����j[�>1�I�$+�S5u+��<�C��6̞�� �!0��:X 0[��=�Q��2�֚��aK񖠨��d�Xi�3ccF���
���e�w����ք��R�C���"F�b��?�9��_�о=��&�;w�(���!�
�Y>k�sZ�s��^��.N��73�J���3�H���T�#V��Q޴��t�<�@Ck�!@D0�N�N������۠��o܈֋/K�Vu�6��o܇ύ�*��� �gqB�����y\�E·���\(�y�-E`��S�?�?��v�&��}ɵ��-zNN����p��M ��^��-[P�w���q�ȋ�@kU�c��������8�O/�=c��hsQ���V�K�r�;!���Μ�O����:�(�Hb���wp-9�7�<����gi]uh���5���g�B��.i:�V�XyiW#r�Ʊ���߁3�����E��}�4����8(U��/�0���N�qG�=b����%����`�ؗ���2�/e�?&�;��4Nu#��6�>���j9�a�<6��YY�w����S���l�����A$��@��%��$V��a��&�b\�j��VC�+9�~�:���L�b����%N�q�qQ�y6?��7�^r1O��@�1��v:jcN�r2�D����X�T�\Mz�y����/�[��2˧�pX�+��|<n,1�<�|��c�u�˳8��a�S��x�mp����i��"j<��Fk{�V�	T�.aQ�`x}	��vc����[�щ�s�E��F�._����p�o�9˽�����֏#"�L|rq؉���U+b㎝�z�}��MA��˄���!����K�;��M��>�FAz3���
:G?��7^��b;�䵋���1s�@�Ӏ�jk��Sｋd��m��u�.��8�������t��;�������Oq�G?�s�Ν;����-&h����m,��S����"���jXG����ո�1�NtK	�;�P@���� �/�S���"Ar�D�*u;=�J�h$�G䱤19������[ᎌ#�0}�V����2�#��?q��N,>E.�Hd�|��P�j��Sy�x���sz���M�#@?{�nl~�Ul`��>�/e,���8����P���v`�9
OB�%&-���ôi3�i��yz�3�%=ߌܖN/1��k�{|KB�I6D%Q?�T\Fד,�-`�}�<-�{�Y���]̅!:CC��}�>�-`���/�x*X�@&!FVxK�옪�L_�3�G��*�@�*�3��;=]��QEb���� �����NE͂���n,�cff�N�5�<��)Tw�D�]��<��¤k	�����p�?r/P,a��.�y�^3_@ʢ=����KNHˣu-��Y�#&f�a�Ta������<f	�K�9[6����ۜcvJU�v䵶Ly!o��ix�*��K��{�"b�v����C�X6O_��=�Q�:K0���CB�.99�<���4ڇ�D��o������4f>9���`x�&�	�oٱg^yW��M�����������Q��t"z�<i��L���H�"!k$RȨ�l���WCA�T��J��7�f�����<2��ut��t�o~�~���ȵ���_�����Q!G��Q��ˑ�>?O�X�P�i��4�����I2�Y|.��(�k������>�/���?�?���q����C�X�����a @\�&mQ�j���{j�Ϝ�Ĺ�^pqȳ�S�ng�4WB�#PՏռ�@� �K��TU�w?!g�v����39�1��O 6!uLa�L�5������9]l¡t]_KU�r�D�H����8bg��T$s��-�F��@�'���J&t1�RQn���)P��%��1/_9�+�����p7n�9>
�\Fa�:�[6c������_'=���������ѵq��GY�4��_|�w�'D��9Ĳ��|�!L�s�8F)9}��v�����ā(�5�/Πu�$�F����=�	\�2ݫ���xK"뢥�{�ȸV^6#1T�}o�_�x	�~�,vn���c�?Ƈ?�ʝ6nܳ[t惓�n�(�C�\r�"E��sCOO��<M*��JȤ&�"D�J	b%q�$����X���p��4DG��K��Ǒ$.��zHn��� ��#R��Z㵁SG�\Z�ONK�ӕ�)��}�<哋(F9s��1�9rn��g����8ēt��#��9	By�X�����>�/4ΝG��9����ѣ���4�F�I,̶m��x��6� �V,�I�,+����m��o���۳|%[Ŋ�R�~�ɾkhY{�J�3�
�j&m�V�<�mj
��4
��Nlv)�Wj���!�zM���9z)[�M^���f�|9�5��������Ϩ�_�����D!X�����T��V�r��h������QT��y;��+==c9(�����#П J�����ظkܴ���y|��#�:<�΍W]��CC6z�A���z�,�����Yr4��w�Z-�.]����H�,B���0��d�n}c0�.�,[�]�)�,N�CN����q��F�>A�v��r:b�YÀ �B��D��/���Ndz\q
(+cL�l|n���D�; #�][s"���0����X���Yݢ?Y �<�]��&�	H�X�vMuѽg��������'���G�X�^_�T$R4�јc����%{�jK�E|��P�g��oϹ�}t���L[�f��X���� }`�f�H ��h�D�Sl_��G
iR+�v���m�aܑ�h��8��� �D�w�f��t5U-�B���t�LyS��H~�|�MJK�E�	�ƒv�����Н�	M�][1��S��J`n���Jˀz��Yc���%{��l2�׳���fi�4�K��C{<(Ň�l��?f!!o��z�/�Ak̽���!FFѠ{2O�Hm���Q��0X;�Nyj�(֍�E2Wj���҃�ED�C�"C��k�yjg^�c,�}�"�� ���F��N����S�4f§�]�ˢ,����y�vCCZ�&��I����1��U�}ξ�6�=n~#M���@�փϻ`�	o<�s�f�_��6�q)b�4��:Y@&kY��|���;�ϕ~���%�o�ԕ���=<��0ta�9Vċi��g8�2t���i8�|q��|v�C�ֺJ�T�Sqv[A��8�����M��{���f�[��MQr��^�M�7�Yz7M��#���;���A���>��>�ϵ���'��<I���$�	bm�f�ȼ�
p{�>`#�M�s�0�,�n�+�edL�u�㌩�Y�Fmb���F��*��X�a�����X��F05������[.�ȖP��]ᰩ�G"Z�,K*�-'�v��
=r�e�b ��O����C`��j?�$1�+�����p� �t]��X������pb�Ll�G��t�az��`�6����%����:Y[�f&��t?8tn�0c�2XƉL��ġ/b:�)j��$��d�2�N���e��й�{	9����<���Ep���k ��2������A E���=��(�M��&��Sƅ�	k�C9��-�:�X���zK-Q�t�92�]��HCz��A��,�?�F
�׏�O�_�׳���A���U��ߏڃ߀�m��!y�m\x�7�.c�#J�Z�X���~=I� :��&��2L)4��>�O��>ת<:��W��is�N߸��[��!.��zY�v��o���Q,'�V!O]UN3+OT�8�Ft�3�vt�,$�YƹY�j�*zL԰�i���}7݌��������D��08H�O.�؛�w�e)s}���1�9#}�(߮�1Wh&����YٔP'��-�O"��/MU�-/��D��q��4��%�ntdĜM��[R�f�t~=v���@�L �%r��S�~YQ�����KZ�,C!ʼwA�T�3@�5p��?��B��kօ���"㐃aD��A`n�;�"`'Q&�qM9"I����W.Y�i�24����*`�o�&��[��`��-S�I�rX�na�Q"bH|l��ӛx ���4�Q�|+l='ce�>�3��DG�]�c�'��М�J
߅����o_���<�kC(�"q�-�*,/����/�_�[ܗޢ���΀��sm ��\��m.\nF�}����Sc���TKU�B����d:�����]U?���-���լpr�W^�6�Y�PU�H�����4�!�J��u+�[ �Ts����p�x�����z�F�+!�kX�W����}Y�ym͟(�q�׿3�q�@��
!Ɋ�x-[�:W��6���ǈms��f�f��X	��!Lу�Fc��V����In�
��r��)��Y��r�r_�}��dC��٩K�]l����g�R��u�~k��}*��3��^����	h��5\j�C~O�>�JG��ڵ�<E��Z�0h+�QU��g��~M�]���@�z����$��Ex`��q$�C�L?��_F*a�+�����ݸ0e:�G�F��q��?Go,���M�?|/��N�h�=��}!����S_[�íð�@��rKH�[��}����}�5�PH7�\!��F7/����y�K`��3ŀ���q^:�HV����,?ij*�)��ܧ�>A�����P?{��*&cp懗Y6r&L��G�{�����X#V��̺Xc<͘�N��[(����YK�J�2f�%�f�(��5�7<�es�#��?T�Òs�O�K��H*���=`k�\%�%��9o�������\Q���B�G.E�Y0��R������I�9Us�Y�Er�,�#�I�q�P�s��,<�mK�\^�����3�F����P-��Becs�`8��k����@���1�?Z欉�|߳�;O����}E�h�uY�_�F�&���!�z��-�ͩih��s��D+"M��ŉ��g@�%��O��/}r����M;��tQ���59�t]��.�	�^F�(������:�Q�i���
��=�`��1����������{���+9L��ފ�GM��T�c�z�[�tIU�.�h�U��(�y��v�k��p�k�<J7��<��qW'�d1�3��
�=�1���al݀ g�Yjڡ�3��.�n��|^�]��X�K�gΡjZ�&jl+��Տ���B%�����y
�+�j�-�|�Ž#U����\P&��D�>��o������2$�|����"]�D��|#����j�����J�XZ�O�&�F��fN�&�qK]k������eBAr@�m]]��eٰ�,�������ZP��6�k��Q�4Qk���S�L%�1<Z߀+�e�K$)
��ǩK���T�щ��l�ģ��I�܂r��������Kȅ�n��/��;MT�s���}�$?�k�%:�b,�,k��wb�����Vm ��=㐞���[GK���Qxϰa�>W�U5�Y��t�9,ip8�6���U�0Q�hZ�7-Sr�, �uzi���@\�Q�@�anو�S����zĎK��%�\ƦJX���G�Ο��Uj2��N�	�(�jYv��ꏰ���6"�J?mХYx8Y�{]&�eC��e^��C��}o][�y��"c�]s?"�g�)�2��S#�8R�H�7�eB?�!2ɧ�#�g"Ks�;!�g*�V����W�Q{[�Lk/uũ��_d���?���K������yr�f톺��:FYpY�ג蓣[ȓ�ҹ:����F�#f}�����9,�r��s�7	�Y=��T�c�8���9V��������w�kM�� �2T���]c�'b`���w�#[\���x�L�)�'�fn���bH�k���d��K��X���;o�\h%}��
�3��\�.EW�|/�^B��Wt�������"�����������KZ����FgU�Yn����\�%���x����~mv��:���DH�X[I§��e?N3T^��T�٤*4�e"wB��5��~ޣ�DA��1_[��`d���0ʲ�A@�'W�kz�JW5�i�t�4ve*z+]���5g�}��uQ��h�iˬ�����V�zu������j��[�5�y�{s�,׵~����U~ސ1��.E*��=�����P g�oyh�����T����r�z��	��&��>�PFw��1�y/��N�w�q�]?�%��\�t6�>��6 �}�j�,88ݎ�d�E�@��x�|�{ĉ�AY+b6�r��Q�R�P�4�!ǁ���+�as���::��e,�ş������1�<��XN�ƽ����i�v�x���2}���sIY���e@l�米��ON�F_��\�i�
~���#[�dNz�1�����t$X^�}���5�,|**�K�޵��\K�'Χ�����ׂ�0���5=�n���7��@��5N\_��.M����4������T����ZP�罯t�*��?�k� �]�5?!�,�ϒ�&ϰgMxi�K������x|��0���E�t�|�+�se�N�wm��G@i����O�9w	yv�;�!��,a$W�_�v�[�si�\�5=l�:����S6x�bg�#9�e�蓞�떁�l'����5'�8�=h2јI��Uh�����,)
��f�I����P��#Ј`[���U�2M��Yyt�M`���ظ���<����Z�¶�@��1�,�ώ:��<��*<Ӑ�1�QY%�� �����~kק~����3C�RE�J������'�k�d�7�KЫ��4��F�N�u���&Ľ�O3�z�a����U��XCe���s�w������.�c��C���QbyO��I2A >|��]�%�k���3�Y�\�RXӾ��y/V#ٯ���k�"cYHu����w��d.�n=��#y�]V�+W��%�~[��t�CNKI��d#�ߍ�-�!���L#�jc�4*�rE��_����e�����CN��aj�U:~ꓓ��_5�3��/� ��b��Y�ė| ��4�k)�;����+�	%TH�ys���9�ܺc�Ff��u�y�&K�2� �f��<ZҶ�l�s��dR_���# ��R`i6�ȡUƶ���[o"d�;�$��g)^5�[m�����Z؁�#��k����کS(�=���`O2V��j�����0������$���y��qe�?z6�·~ DRSH����NW�g�ni�C/�ZW�ݓmɽgs�3�f��������}�gy�~.�S4YT���5E ���=������3�.�#{A�J*��_��[9Ɗ_���S!�t5�����Av-=S��OS�/Y�/�z�@�y:��ۂ燘o,�1���8�i����7�ݿF��<&�n���s���|TY���N�S)�{�7�����X�c�h!��W�>��W_��6 �]��}�)�	�i[O����oG,w����"��q���(�Ҽ!���El����<n� 4败'Zw\�ʴ��,'13�@�y�6'�8&n�x�1�T3��kH����#�>���#(�t�����:ofq�����6����"�A��S8��g0�ʫ�"Th�-�g9Q�"N����¬%��>��_-��?T5�:����_���Z Ҕ"������p�Yk(h�iJ�Rь���%�3A��a��*��~^[�G³Z�d�'����:R ����YHdb�Z�ǲ4U�f�R8#��s���𹜭�����)H����o�Ѥ�y�iv�k��2��~U��gdz����Y4������f!֔$�U��k�Ī�%y�D�0�D��!g��cg�󞆩-ף|�cj����F��u��/���>��7h���#_���dlj�U������=:�3a��C�P�u;v�������m �s�j�.E�y!��?OL{��Q�Z��cL��}�`�,Hf�'�s�yr��R�i�>�`�K�X�h."��y����y�6��W�S
�x���0�0G 1z� *��-�f d��$��w�?��aP�B�V��ν�[ӗ���S��9��k@xM1hp��}�_���p�+�=}V��q�ג��a�bg���m]�|���?�*I�X�n5t��9K#K���((����I�/�Y�]��d-.b�M��\s��K�}ח���}���{���r� Q�|2 Q#Vy��A���=r�G��(�.Ĵ��,�����,��"'t�+fLrxu#F��D��a��/:��|�H�MP����mV�}���?r�����g 	;0��S00,�����{!�t����[�����J>1*[��J�T�'!M:�"Շ�����_v�W����+W) !$D�� �m������;����f��wf��q:�;�n�n����`0Ƙ,�P�*W�����~���)!a�}ۖT�]T��/�����gCӬ9����T��1��`Հۨ����(��YYG���p��0����/`��gє���pN�8�6�9�db���k��Y�)�H�2�ձ�K��A4�?��e���q��Y\�� �A%��g�'U��l�*��h�\�B>������3�����>��^K�8{�"���k�)��L�vz�TwN`�AV��O��"���F�8�F'{�|/�2:wp�[|�������u�*�{c?W�xj�ԢH�g��--!�D�������M���x����l�����ϟ��#�/����4��*�n��D����<߽xl=��b</��]��"-����l1�/��[K�p �'e�Q��$�w��I	�C�`]N�"��V�KSێ�{f�1w��4�Z$hE��>Š��%*	���殈��w���5�b烟��A�ScM�|�=,;�+8#��hڣ���cP�`��P���Y7�@��m�D���(g�0��ie���]���Sh.�`�Q��]��K�6E�l.�VY�&���?x}�6���K����l*��
q���g�}O�_�:�i��D��x��Imqd��ʹ�;LŔ@lp=��Q(S���(yrC�9}��s�G9+����<x��w���X��p���U��ZKG�<y~��i���cx����s�$*�r-&ĹIB�}�S�?}�w���o|ӝuD���|�V��o=+np�\���l����f���彶 �2_�>�"z��Y�Y|['I�0W�O�:]�Ij�0=�a,~YJw��A�Z3�9�������A�%�� @�:>����s߽���>xSsb��(jbo����K�Uy�TV��u�xv�w�vZ%7]�15�[Bed�?�tP���	,��G8��crq	�-����ܥb8�t��!���:����)�Opl��#2�ύ�?�f�ݫ��fP���;�{<Hc����9�t�꿻8oxNF9S��$@��J̞�m9��CZ�-(�wPF�q������٬���@���Yk*�B��8�I�Ǡݑ#L����&m�Ou�$�w����'��1���+�8B�䄈3�vhʅI�d7K�E�O�y]���u��x��=���g��.ϵ��z����C�*�;����\?�y�A�ي�G���ۜ���Hk��i��X3g�ܡ����ň�P.�އ�>,�}/�+� �_���~lB^.qF���g?��_���b{PU��@���FU#��M7�%/̄6d;�К/�]����q��η����aV�=]$�m�ӓV������������7&��V9g�sg�_7�nmS/���L�sr*
�0����\1�Nrea%V�R	�|>DQr�9���q8߉l��P��o��9�A=�GRG9 'K8f��v?_�T�{-
�'�O�X ��6fr�\��x;��m���x��_�kLJ�_����l�vg�*� źl3��hN��}z��u�;����i��"�U��[��w���ֺ���_�kB��/9�Q�������E�@-�N�m��)v��i\b���������Λg1.�?BK����ǉ0��D��}�+p�\#���Q0��;�w3��*�]{^=�'N��=��cPm`�9�ѹ�{7&XOtm���q��GӜ��ı������Tg�Db���Ѱ�b܎�w��ؤmN�P&�"�����~ؿ����/RR8-��9�\;S��1F�%
����+�ch$[�ϑ���-{�&ˇ�/����]z�{���weE8f>�~�}|��-��1��b�L�V8���}�<�42乸�
��_I��!�v�Y
L��Ήz��@��kS8sޭ#)<���������^�T�wQ���N�<р�|F~J�iW��1�nMo+�~��-@���S1��D���y��34)�~3��P���j�(\#�ܵQY��n���u�j�wŸ������ƾ;n�̽���+�su���EW�W����8R&=jM��~���+X�_G#��,gx�x ̓ש՚��kX����d=3=}���_����؞ǘ#�=�`���f�°�I�������P|E_�����,��$�9�=����t�H�댐�L�Z����N� d�j��{�� �[ֲm�\u�]�j}�Z�VMIǦև�qk��|���I��x� <*.3RWWy�����KǁNC����t=�S��4;e_u� ����ߣP'�O��"ա8	�s��T�I�?٨#���KE���=��ڏ�9��'h�Mt�k����p167��m~."w1u�N��|_�#]��t�{�m�?����t-<������;yv�*����V+v�4,�i#�j���(���l��be`�6�5��*D_x� z1=���@,ۣ>����r���:��kTٷ3�܊��<��R�Z������.g��_Z.��g}3����������1�����J�k�6uL��K�CY:��*��6�t)�`���ޔ�.AV���z�������zF<����gA��O�2X�7P�U͘�T@8K6�d����?�){�͎�=��˰\�mK� ;bkd���|/���N���[tL�?w���+E�Q�f �}a()���r<�*��^*ġ� i#������ESB�.�Ž����/��8���OT���1V	������[8�ϩוm���z���_�
[��Z[�~�w?�Y��]t�D�R��f�_���=n�Ù�F��gHw7I�k��5Q���2���� ������$�h¹V��*,!�F����%E�n���
�F0;��{���7�b~u7�~��^���2  ��IDAT�L�_Py��%���w�d<FRqK?�>����D�k���%�:���2+J+�j�夲MZ��r��b]�(0l5������7��өcj���k!�=�7r+���XG��Fa��^$_��跺��(���	f%Hä�˹��%��<g��0��tVy`��t�G	����8!З���H��JEA���ڶF�@�=�T9�qdXS�=�bs��#Yi���tߍ���wb��g��vOm�M�@�����D�+S�fU�)��M�8p��Ef�o�3ڊy�r�ޖi���]�פDi���*i�w���ܷ#��$��f4^8r�EaAo�ۤ5!)��Z*�`j��ǎa��Y�/���[?���Cp��22� ]�~'��(p1P��q�A��w7N��
����5_�V�T���ׅ_�GXb���跾�����$��)]ӌJr���j��j��9Nyҹ�|�Ujk}�R�SW�n�N�w�Z3��;X�	CK2�a@.%#Y����kw�@O}���
���7�2+��t�F�kU�����԰u L�{�8��C�.��3��[�29��Z����W��Ь7����t��Ε��ewǬj&@聂� <���c�EU'B]~r#|�u�X=�wm�o�c7݂����~�X���ɺ�_��V�Q����OL�wdw��2u���g�۟�b�_Nk�/�u�5:�
p�I�H԰��9_����E�$N�b��P��֕M��ٔ��~`1�8�A���F��ӭ��9�SG�b��<���"�[n@8;��&��3�@�Q6R��ױ��`�����}P���HD#�@4V����`�������ha�C�NK�� ��J�
��
�x��Ρx�%���f-��ȥ�r��Qz���CY��U)-Ј���v�mU�@3*��A"�9!W���]�^n����.U���s�C�}Q���f����Mxvn{nHm���^��ѽS�C�#��F�a�Z���� P@��Y`?=�%�3�gj������!����'��NrQ"����-�㋘Z0�'��e��K�5��}8�������JU�u��j�]3�O8E��l~����JԾu�]8��-��岶 �2[�U�%bʲ^�	���2��K�9ӏ)\�����ۦ��t!0�ϝ��'9�oV���˯��U����NK�U]:��C��߻��"�J��T4�:�cs�
*{�D�5�ӳ~��J�v�Ħ�Ι��:N~����0.�&=9��Lc�0�Ď�	�x:�k�I����p�܀ԝ?�}�)6Z*({���z馟7ް��d�[C@�@I\�	���QXA=�!�}��?���Ԉ��$�Q�H���74⵵��z9�4b��|�K"|I`���M����T���/��m{e��
�p�yO �)�0Q�׵Ʈ@����gS�7����᳎��K ��f���q��.'�}�8Z/���C��1�>4t�|�oƻO���"�] S!�-�k=LVk��v��� O^�V:������u��-@����G�-�y�f� ��N<x��d;f���|�^n'��cDa[�l�$1�g��#�I���sH�^u|��xU�u�o�����E�֋�����n;$H[�(]5�RW�\FS�t=�B��ֻ:��p�gܽ#���S߄��4����Pi�CAX�Y���!'��oF�Y@�mx><{�Q4힝�h���|����/8���O���#g��r@���CJ��zg8`��N����4O���s;�dāд���Y^5R�M�y.�~��c#��kH;}=���Uy��)Me;좨��[<��%�(��?��1M�<;>e�I7�]���aU���{�ˈ���W��[�=�Zsgz�?[1��q40�7������h��|Tj5��Zʞϕ���g#sMi�:+�c�Fr<W�_�I/N����p�N�Y�)�cO���~^����>����w?@JM�:��6���Y�k27�y��9�n���\���;�R�����h��$@.�Ntw��A��w�YTK{:�3qM��C9Ak�r;fT'�h��	�<31�5��5�4�Ԓ}�b���PeW;�~�,�*��� ��� x�A*F/P�r���b�d,�ِ�vyo���!?��z*r�pY`�$�/�z��ߑ�˔`��*��H��sF����k�.�S����[c�(ѬTvq�z��(�!�1:􆎊c����������(��|����WvDX��-y�zq��	����]L��gN!�{��"U�KX�f�]"˚ :�L���$9��=�!o���s�;�^��t�sP�GI�l �:|�^����}0��`�5~�O4
��S��ʊN��D�����>�P��My]S��S�r��U�^yK�6Nʅ{�����u|�;0wϧQ�1��?�!��;��؃���k�`���)ׯ�w��֟�s��Ѝ	���[f�rY[w�2Y��K�-9�S��ƕ4���;�+����'�F�cc؈D����a��Ig���+GԨb��8#�G���p�����7ې�Ո<�dh���֙�ĘVe��@��G�W/b�׿���$�!.y>���d|����Y�	It�	ټ��]�iw��ӎ���L���������(�Qb��s���r&_��9���|��!���a�~�LY�L3���V��Ud��u�����}+aEG���j��W�ߓ\�QS�uwN�c�Ek��aӟw��G/�<������Z&b�;�lC>�#ϣ���$&��2�v�,�	r��7��c�?�k����!X77DS�������{�C���ӯ���X{n8�=��n�N(�i�C��X��o������W�q�ı(��]q�����{�+���e�� �4�u��C������K}m�e�B��R#��d�dZ�J|q˄�f����|�<�/Kp�>�ڈG#%��GU~O��W��yg��`�u
���gv����ŀ���h��u�h̰����8���a�D�1XM�]h ��+Y��I��� ۔2S"H}y�l��D����l� ��>�A-צ��O�L��4xFF����h��,9+aіQ4�uK����+�yC��W��5�Ἣ0܇<5:�w��c�Vd�d���ݖ�,i��$Ν9���o������DS�t(U��#���\��QnS�c)e{��Or7t�9�{��rGx�<�~�[�(0C`g���ýN�����$���U%��觱���cEm��A/x��g��S�ZU�~��ݘ��_{vc��B��q�;g1}ݍ����TG�fU��I����}b"<��x(p��<�}_6�S�F�����w9�-@�ֱG� �.k�y�9Yz�J��t�>1M5�v���I�+�]76C/��\aIiC�5�R#Z�!�����UL(�~�U�tV0W�1~���b�_dCHN�L����8����o���P'X�]���y&�j�a1�XW�\�O���`R�(�5ۤ^�D�3tL���^ym����C97=GR�8�, }c	dNYY0��e����׶���Vƫv�J^����AA:�ɦ�*�������ct�jͺ���-�vO�ݵ'<Ϭƺ�te�^Iqv���B�O�W9��p3#�&�}f�|~鬸՚iE[K�9汑d��_��Ԩ���&����ݞj��T���"���)�����|��s��.#�tΜ�����`3�܈m�=�P�yuI�+� G��>��
j�7�M������ew/�>s�A6�sg�o�Kqm�e��bdZ�6zi��jC���y^\;��n%O5��5�#��`�M����<^�]M���zk�q��4*�8r,!뎎�{�u1�8{�8^�ǿ��b�w|�b�S���� /6�a��I������y�#��}�h"9܁��qf�c�ƙr�2�J	�n"���lXnk�&H-��L��;�p ����׌����˹�b��z�a�ad��#���9� 7�ޅI�;�֛+`9p�)�2�/p0eݚ)sq��Mīk���;�Q�"�c����z���ŒL�>�|��1�5%ת��H�q6�h]g�5�z�s*/;&
��+A�4� �9�%E"�cO} ��v���"DՊ{���:3���c{g�3r���'7�Ⱦ֏A���:�Nw1������i�Aw	�j�8�k\$��`}a�A�=��oq��a9���~v��������/��ֺt��_����}�����i�Ź�R��m101��#i$jLa��<f�5�������<�"KH�����5�`T	e����5�����U��/��ڣ\���t0��ϰ�c�*�%��7�p�9Ӊ	Q�A�QI���׸p�y9yh�>��,o�K��ʏv�Wj���A�O��{y�}���U�W<S�!$��A�b�����cqKu�m��2���	�#��|�S�*�"��Qo
��0G��ة<�k�J��U�� �9Ɩ�_JĔ7�9G�"��S��h73)}�fGFK���Gs��$��G������� 6� �zC����3�s���XS��3�q��;��D�/͍�M�{�V*��Q�5B�b�^�S��YL�_�󺖏Z�x�=/�1.q#,�#����%p�.ײ�`:�V���Ӂ��rܿ�ڎ�oB���w݃��m1�/յ��:���uPCO"W�r<dkY��v���]���o�j�T�0�P�gKB�f�������5sLu�9Y�fb�:9��L��H�q���D8�"����5��x��9�s�<O@i�o��ŧ���|�j���r�M9�)y�����V��D���^�W8
�@��)�B�'�1T���NK���H��d}M�[ F���β�C��s����j|">݅�w���H</0A�n�{��XX?�ʎ�N S�d�sh�\⤙1D{�T���F���  S�-����(.�Zr��0��~����##�ʄ aπ')�<���c�FP�������<��{dQF_1����s3=о���U��,OT�h*����
��đ!��/:,A�Z�g>�k!�Mǹ/�(�~��Θ\	���r]*.[�(u,wP��.����8x�v�g~DQ�%��PY_���Cud���g��o���+r2��P����ֺt��_�kRI& ��4��<�T��mo6*�������)͓���}�|4b�XA}nؖ��(�uģX���?U�GAJ��v�/1v�P����&�nR���Q��u��A����A�k��?�3�'�b6����� ���u���ژ��V	A����ZC��ƤD,�|���q:�G�@(8r�U���1&����Q|���dX�Xel����w)1L�X�'����~�߈�e-���L��L�'�����y�r=]�k�+A˴�YU@���_ņ�c��u����.׻�s٧:�+jG���s�Q_=4�/6�S2�/D����J���r�ܬf����b�9PG�ז3{!7 r#-�佞ћ�r-!��؎�g�V�*���̘ܳВ�7���9��\ff ,��ƑTǰ�'=x�fb����2��	������8PՆ ������T�>�oq&���(��ɏ�qTd�'$Jߵ�_�k�/��ƣ�$k�0�7˶���I���6��F�Q`si��c���F��ǜIb�i-2�jW1�ku���0����r':b̼��1C����*���"{�Et�z�Z���6����5`׵(:��^y;�S+��"����GQ=x�ѣ8����pb^�ĵ�o�����=}K�zZ�����s�AL<�l����Kc��}�m,��E�:�C1̃Bg����J2�?S@�cK�Z��	��W�`�^����8f�Th���Rm3�@2��˵�* �y+0)��M�Q�7��ퟃ��.?��?�y ��&������QNs��JI�f��&2������:�����}�!.�Fh��
�Vq�u7��؃1~H�·�W��"���a5�|I����lbbrJ9��N�/�h�7@�~Bj/P�X'ҹ��y��0@���+vÿ�`�nt����;�1}�N�����[G��@�?�K<�%N'˯n:�㲭W��[I�Ρ9�p��~��-@�D�T"�ȋW10�X�{����x!+%R5�M�1J�$�K�XHdk��F��䴞|��ݏm���{��.AU,*��U��*�m03�S+K�%}LJ䜴����ɿ���1���c(�D�IŰ��n�X}�y�N. �*ؿ�Zx�߁��i�����2>�[���n�0�;�|3={��5��<�[���ֈy$�I3�3]�s�rM�&:�g���L��ۯ�?1����	J����*�_{��ä��:�!�0�r�vB0u\�H�P�%�7��0o�.#��	ԔL��"��B�L������f����}���K��& �vǥ�4C��Qg���%� ���EX2����F��jj>�����I"ci�}k��%1I��wPU<%&�F�©mW�75�N�#�2D���8����94��	P�z���Tn��$mLVj�n��7�;���q3�.%�����/��ui�-@�ב'��jh=�fg���e�YZ���n4��A�%A��ڠs�_�Fk��Α
5�`�08|�ڄ���5�FU���WqR"��n�4�n�~����Oc��wpt�,�� �4��p��ʈ�*8��K���>���16d�u���H�?�H4X0|z�		[X��* u�m�A��z$cx���������{p��3�0{���?���cj�=�-]��8p�L#��Ss8-Q`�c�n���"�� ���*��>F	�+���.b��Wp��g���[b�sT�?M���\k�·��ٵ��]l���q�L�F"�Ds[�_���t�&ãZ #D;���I�uF�o�r:�{����{��8T%��ķ�h�\��ij��F���w{(uݫ�>��~��VL=���9���k׉\˴�A*����t��Z��.p`�^uũ�pW���{��*�����Y�I�w�]�`��{ޔ�_��SOnm�ۊ�/ŵ�࢈D���\��Y-K����.*M�k'bZ�!��&�֑���-�|���cX�܂�[����*�J�k���H�2�=|���uT:u�n����k�[T� o�y㵸�+_�����>8��?�!N>�K,,���O�o��c'<����:a���B>.�Ҡ	o�vt�1�>�d����QA����x��?����$J�w��(�l���Ze�av����=jy.>��\��f\���Q��3���Գ~��M+[�>��s��X��&�����wb��?��O�g���TA� +��&r,���-��^����FA+�2����kz���avx�~o������GU�\ʹ�g����u(��^|��ץr��iŋ���a��+`W��٪'F�!�RfB8��_r�'��������]	ȴD����u�c����-��h���u����w�z�X~����F�F�����D��5��s����j����$�%��)qXq�Q��oE����Kl���c�%�j�/u�,���%_�8�ܶJ�ںة Y" �r�g)q����K=۪�l6�0�Ι>g�d��蛙�4����dR5�9ﺊbj���G��߁��48����{�(^��ߠ��z\���7���"^O��ʛ���_��v����~X������������J J'f�IS���\"mG����_�_�۸�z�����^������������c��9����vv^Ȱ���Jg�3��yT�ef�k�Yя��|��5)j�����-��*�	��и��y�!W_m��cyO�.�K��9�;7��}����ȾXz�_����4�_����]�u��g��`6����D��n�m���;v�_�6"�{�ƕ�m��n�1�ߘ�6�?׿,������f~����jPW��	z�<��YH��+u2�w��FB\JYW�WU�J%0�<�!K5r���ן���\϶�-g0�����1���v��s��B�Ibq8Y�^�3.��b����ʚ��Y�����3��c���R�:P)t�(Ĺ�ʦ��������Y�d�u^�Ku��7��D��
m�?ǵ�ؚ�B���S�5/�n�|Q�gvת�� 0�D�	`v
��>�N�ᱠWC7�!��w�z)M�o��%����<V�kG�=����c#{�w5�pQ&A��	��,'�����N����g�ڿ�;�ً����!��A��j���ȫ@�QMh�P>C�e����h��`�>�h�^��?�_=�m�^���I�YS�����t3|�O��գ�Q�9Q���k4��F�F�ض%#���&�T�X��Q��n�/��cL����:C��L��:aG��}��� ���gl�p��Nr�I�X em�5�<uT;c�����P�"�w܂�&�xm��0��QT��+@�w�֑L'��	4[bN-:v���)M><_{�<G�|v���a�p�؝��n���%�n��]�Z���ukt�|��Ua�v7F_�_r?H��3��Y�v�B\̲I��a��7Y��n��T��Z����<��ZCC0��qr$A�Ù	�l7���`�";�1��V�	��g"�cgT��'��/�.�k�����&��[���R�u^I0Ռ��Ǡ� ��dT��ױ-������fQ�wy�U8N�Y9�|L���Kkm�%���Փ
4��q�%����OV=�Q�����^�e2��sg�f��Fr����ߕ��v�t�t�[�W2�O��D7��N�!*u_ga'�6�*�DQ�N�d��cX��ͺ��L�c��x���t�j3C������S^;�R��y�SLG@���`=#wp��8}�^}�U��1��.\u���&+�wa��_c��Q4%*��f~�ƾ�m��#�/��p1��Pm
.&�v����ۅz������W8����]�>��:��P"�����cp���<��4;EΤ��}����h�+᱔�S� �_�՚��^��_�">8�XZ\UQ�Jm��)UF���9�n�HI`���us��<�sR�N��4@aWάG�8����lʴ����33�]U�D����VH��,v�9�#t��U~��Ć���1,0�^.N�?���l)��Ù3���v����ͦ8�t�ƌn��B�}�H����f���GG �W�ŕ7~
�������C�,�&��ғ�W5��s�hf�z�e4�`g�8_��9�Sԥ��}o��r��{���-�Kam�%�t ���iBB�S�{��9f���8����2���Za��Љ?��=ι��d�Ta��!�ɠ#QEG�vZx��G6X�}���C�ʝ�v�mx��/��]��ib�ܱ*��
zu�$b�0�!�
�N��*1��V^?�䧯���Ѯ4��/Шȶ� ���0s�ع��_<��=�Kd�W���U�PմgF��J�"�0�9�c��I�:�ex�
��yQ��H ג� �"�M��M!o�LŅ}(��Y`��Y�9����_�Sr�$��\��c�إ�lFcި�QC\gm3M���r^�Vי��SЌBY�ca!���w�},|��bz�d�ڵ)�mR�ô�y�B�p���ٺ,���Jt�k�	�3`b:�"tU����^$��g�����sĒ�
�f�
q<3���kN͟���:�ھ��qm�OL"j�����5v� %����|_#��0Z<'3�ŕ	��y!�:�W�E�_@���O/#]Z�r'SG����s�/�x�\��q�,`[��G�<��Z:K��m�W�d�֝�D։�|I�z/������▥,�/S���^b!%.�Ơ���6U �)Ώ__�1���1}�.ۿ���bX[BU����2^�'8���(U0s��s�A�t�E���h�|=nx�~��x��TV�$
_Ď�äW��_G����N[Y���{�'ug]����� ���1�tQ۳wL=�+o=O������߾����&���>X늡f�_f"�k���XO&���Z�"��o^[d��zS�W	��]�ݵ�4�빂�˚���y�yX�B�W��y�3h�q'��.�jW��ӭ�g�}��}kvk�f���P`Ɖ�:stl=��1�O�}�V�r &����Ԣ�)�hN��%}�F�!�`�g�|\��(��WhO�D��: �0c����~y^�v�#��Y����������&1�S�N���J�MBe_I�#��Q�Z�@ ��C{~�^Wǚ2E���$ʮ�T"�_K�d���F�-��zz0U��yw��H��˱��͚���y�:=Ԙi(b�M5P�.���|z�-�����q�0֕��c>s�>l�J�_�k�/��ړ��
u�)?)�L��O�)��$iV�	o��L���C�2����66uh>�a��K����4�Z�q��<G�.16���~�G�>=��޽p�{���ɏ�����1X~5�YӅ�ί�G���|���Q�@ �|қB�0��#[_A1pP����0���=����3	0��C�g���T���?�?��'Έ�K��XB,Qy&���c�2�eڝ������3k���^jWA��ՀwK�3׵0������SP��:�i=�y�H � �X��z�A�}�~8��U<JE3�,3L�|�#�g�t��� 6�"gj�Y���)�W����?�����^:�}�5�M�|����=�s"t���I�g�\3����B��|�̙��\L������N֚ kC�y�c���;g���aC��x���y�i�a[sB5�9���k��e��Y J�&��VB��e{�{�hk����XC����`u�{XJR��6�x�^��&q|�0h�b����s�@M�q��፹qtVP�Bo)�?Uuܿ�?)�\%9.N\e�o��m�%�&h,��'d��i�d�-�I��I�1�9����Ӳv�	:��O�vwa$<x$��uql��8��o �&|ΐ^����2������� �THd�l��//��o���W7�&�:Xfyy��>�.Q�m	���vV�� �]T���Gq����"�"`_"��Y�f~�N>	�P�]U����L��@��q9�P"��A[ R�Y��#Ҟ��ԙ��~<���1�F���kn	_��8��囂�a�W	��F�kr�~$d~���3VŞ��E(P!�CԊ�,q��.��=��B3����K�t8x�=����h�
�y��� ���nG��p�G��/l �{:l�pk��&ű�+��7޲�]�!:��H*XF�Uj֝'������2�1�*;`�Y��k��q`J
�_=t8�=V��oRp�Z�1���	�Xgdl��`O"s*�MML���5�d`��S�DVD:������81�4�ϑܡ^,ۯ��c�̻�L60{�����O�۹[�(
0�'ּ.~�[��.��+���D3g|��{h��C��WdhPMr\l��=�cck]�k�/���F�,�?H��M�yr�؀kvD�W�w4}�Uؾj��k �j�-WvH�m�e��є$��Ј�P/<"��D���^��/F(5N~*��{��w$*̍$�D+3�g��.&��E.zr�����8B.��?�B�,ѩD�͞*G��� g�IXXP�,�g�}J��zX}��)A��0K���!���p>u���@#����]0��0�s�)���
b�����$��V7ͼ� ۈT�(��#�F��^��:SN�������������0
Py��Ǝ�>���n�u$NN�ɽ�5*gF@k��}��֥#��J��Z�-�p�wU�����@��b���a�װv򄀓 ��j)��B)�B�u��L󒩿�6�>zK�t����]w�UEI�+��9�:��g����i�K��yӣyγ;J�K� �Q�f�L�J�$!.ё�����q�{+O�u*Rq��r���\����|ѹ�4�q�>O��r����4���zl�Q�F���>.����I��biE^���L���rǦ��\1�gN`��2��5�W]��=���#�a��alj�� L������$�?��ێ�/&��=��~n��ym�E�(�J�ڗ�A��e��G^>�w�̤+ʭQE��]�ldG�h皺-�QֈH����Lt���W�^RnL�2��ܡ�
����P��rL��[QX#��E��؈]9�,������Ԯjl2&�M��h�0�:��_el%���L�,�FTWK�Zg;��y�D3�^Ҹ-L�"��,ƚc�v�Ř3�J��	1�)�햦NcN��{��s��v����J��!F�Cg�΍��j�l+)���JG���V�m�p����ރ\� I��){���
w�;M	�P��0��q�lb�/r6��}����~�>l����������[`�x�uqg㦗Sڜ�\Y���9e�f+X�q\��S�=�����|�<�@��k��� ��U��#�\>;�����Zf�����'�����3SSZ�B��g����>Y.a]�;��;�t�
���P��ǫ����l1��SI'��j����
st�Z]��D6֕k�y�y��Ä*��F�>��~��3�_����O]��>��¥y��И�"q[��[��5'���'f��Y��?�7mqX���D�[Q�E�� �"^�~�1��(b	/Mw�����;�3
=�iRK�!�M)Z�Tb�Z� ��	FK�)k�Ku�2J����G��Za�^r�4x$w�k�;k�Zo�M��ч�����,�̕'�XO}gX*�-ݦ����h(}��>�;8p&�Y�f�T �@�Z�8��X�3��H}3���hV�	��0	|;�p�bl+g��h�����'�}f��� 7l�c����� dI��(��_o`Y���� �n��4��$H��a��N��q	�rͻ�kf���1P����4v�aH� 7�o60�Y��_x+��4���D3>�P9W����=Ǧ!.���׋a:�OF�A�9a鈢H�C�pj��VbU��m�oi������]�$��jcl��ym�mN�t��˅&q���*�`'�t �2��U��X�B��)z>���bg���l�=a�G������D��ZFnV��l}�3o�!�3�a��?@'顺�B)�~�H�y���ko���5w~�ioR�?@��äWG7Y�C�%��d��W�,�;C�]7�Pg�~k]�k�/�5�a%���*�'�j%٣NVkJh�I�ɔ:_2��L����Jc��Z#fO���v����K����#��V��͗���.笛�����P�R��~��)�z?��^ �I2S�'w�͇s��a$�l_.2�z��� ����t��)��8E=zE�ã�ϱ.@�Z��pk;�Dpg�1�c&gf�^_CM��R��J��81S���jrQ�8F�V���m�BY�p(HD����6���;���<�$��9�̈́�ېY�a%3��bFxڔ 
�k՚���Љ��Eu�5ua/w���$��;�	�܃�{�ű3�P���iv��ɮg��n�;L�+k"S3��kh�yyMx��H(��U�af����,���|�ԡ�}��<�*�}�:�Omq��^���a���OpV{*�F�I��p��=�=�/UL��z��jw`V:5�]l���Y3��3���l�Y���	���M.��e!��%#��L?Z���z^�o�_z3�`z�5���������K4g�J���v[�IK�*��	9�f���~��݁�y^ G���������t1:gq�ק�w�,�"I�/�9��m�����D;�F��&b�����v2��i|��f��0�Y�N�y�p?D).���<k8��:��J�Q	�ƪ�׻&:*t@�~�Jcq:R�F����a ����I2��`���[�l|�?��y��iYGS�f{����]�Q���o�Ā&�);�8��mcb�\s���4������S�ͨ�5K��:'B��▗M���5�
f!���N���{Sw~F����.�c���)5�s��R]���eN|m����_?�F�����#�}R5.E�9��8����l�����w��?���'��+�=M�+�QלϏ�N	�F�F��d��g�f
U�P�e�C�Ca|W�������3�)��v3�41f�{n[�<g�l�1e�y��zM��tN�>)�Cu���Zyd:.��9����>|O�I�ת����a'���f\��]���Jb*���s��&�Ό�>Ś��=��%��Ϲ�r�3�<�;������{���Bm:�����[0^k��O~���ql��Q�xj��3����F{:)����!��%�u���ںs��k�u7����/����ۮ
B��g}����Ud���L��ur��k���ӞR�ח�f����tu�DI⺰�,��6S�\��vJ}�kt4��(��I9�#҈xqmI�u���#�iq��=��t+n��A�s���8�l��M�H��'��I<3	�Ѻ�if1�q���r�aa,	�,|M�{i&����4��0*��'���F�2���C�!�w��ֵ̊�A�~XC]g�� W���j�n8�m���,��Z	��td�e�;z�s+�J�$����y%?�駾����Ǿ}W�o���W< Q^���r��1����0�e���M�Ǯ�u�X:�zkk��*NÚ�� ����#���1�ƻ��s����D�0�0�s�ulo�|')����Ѩ�U1#�r�q�)��5�u�Y%lbllg������f
(��=O��4�U��O��-�h��ʇs�-9��5��gK��(��X�3��}����c�_yD&C��v���|nܓg���X�8h�y<� �}{H&��k�p�{?��s/ $�M��N4�9���Å��gw��!9�o{�x���b�0��ϰ�.����z�ˏ+�Ѱ��L�����l��l��d�F��e
QT|$��*D-��Y*��b��n�V�~���$���FJ�0i΀z֌<�'m��:��u	��,פC7��Lx���I�k}4Б�ۭ�4���ވ��B������"ߤR�ߵ�k�,��ʁ٘� �9�H����1b��u� ���u�?��.\ɑ�d33��z9��*Ƒ��Y{�[�6ǵZ��F��1Ly=�E���C�L"�uP�GPG89��{�Es�>���S^��h�NfC�Tݘy:k
�&S@`$�*�q��������Ϝ��-�#uh���f��t3=���{9&�ɱױ��s����������e������v��f:Y�-`.�ǲ��ܑE�.�k��D�tP��gЌ��E�ӭ�8�<��9�M��&&�U"ă�l�S���:^6ߠ���Ψ=PΉ����Pq� x�8r���F������A�RU���/L���};��
KOv��.`����%�h�5��ف�;o@p�~,�s���ƕ�_��n���,>���c␭��!�Nj��k��_7�����'Ǧ-rC�����[���jm�E�*!l@W�5��Yq�\���9A+�%�ÿڬ"�1���$���z�iWu���
���H1�� �Ӊ1�.@�NŨ*��h�m6j�-I�FF�T)��Dۦ=�L����̳oZ�L�{�ƍF��(w��9�lv@�80�HC�Xyo��܆��U*��[�\�cm�Ύm�*��l�%w��UV��cB���ǆ���I	�w>ǉjjۀ	L�?�4�6Qyư�gmKc͟�>���̵��B��{6�֋��v�T��E� =�ɤ��;���@>5��7��K��]��3��yt <3@$#�ε���;��8x~��i\}�ض{s�{6��Z�on]�m��<�Օ_T�-ٹ����c�/�c�W���Q�t�K9
l��2v���I��5#��~	����F�@��J]e�=yV��7/�,C�tj��V7O��TS�T�]%�j�_=¡ק�Vv9��������1 ��`�lAP�� RF�
�#fH�,�3�y�q>�6�����퀚.1e=��i�u�#t2��=�c��#L�E#w��}f�n�n����3O�	'u����}!�J ����������������ۿ�[���U;~
�^��Z���7��^7+O�����u�n�3Yݚ�~ѭ-@��֑�<����$���yq`u?9�hn��'N��
L�cU^4��0u���yõݥb2�&]��."�Θ� t��C���dq�JK�#ۺ:�������:Ԃ��X�մ����b3�ʊ˻%���Φ��oT��!i&�ў�����ϳ��2}9�ÇB1wh�G~c�r�Y(K&m�����Z�5��HC�x��;yy�/�-��9�1�u�/v��d�F�/�`���5J}qx|�$B�������3O'���\S�S�~�d;��K��c������>kڥ�<y��S������3��-3��Z�}���#ؾs'&�f�s�N9�LY��%/*��*�g/��7���*���o��������ԕ͵%��ef�����>��%ʹ����~��׃�Ʊ��J�(��eo���\3JTZ�����򲊰Щ� �'���$F9s�|,J�6yl����lM��$G�5|��;�u ���^WG���A0:%��@��\��7z�s��p̮���S�*��󒨣fv�ھ}�~��7yFUR�b�.�c����9:��q��{��>��4�a�8��J�'����\�WH�m�}�����=�c�V�E�� �"[�|�9b����	�|����o�� � �5p4�HcrW�Q�ί�����3X�H��E?�a�z=TkL�nGon��N���k�W{��� ��)BHb<u��4*����Z *�!~�fV3�!�34�&���[����z'���<�(y�*r��<ߴi����d
nPH���</�;ڛN�%��%��V\��t�t,�P[��/�-!�R�܏���1>z��� �*JP��3�f ���RB�ɂ86�cT!��>;�[�W���H�(�7X�e�\�IY!)�:{�����x��_c��B �C��i����&�a�&m���i4Nv��vp@�F�r,�C%� ��r�&��l���:*����=���:*�C`c-�5���� k)?�DŲ5Ӕ)Xj����c8#��&��<�y�����T�U^�c8&0����(�%}8�RX����k=�!eāV�~�c�@"jɩH�|�M7���ϕ A@���a�u�|�¢8�c��5sU9����;����E��
�Ge�d���,'��V�~Q�-@���_������Ê���ц�6��|�`W���_@��;q��t��ލ��u[XC/˱�`r\��JdJabc���*ҥU�O-�!h��*��$�R��;l���8^�#*[��*mX>2�CD
#b�� ���{5��wa6�懲~��t-�a�u���AO�� n���)M/��X+um�N��?��6���V�)#V�>�lh� /9�)[��85�'}���_�d�M�ƥA��p���J�sa�FN�){�h33�㬆����zy�,�j�9�3_֎����h�>�~��}��:�����9Y�e��9��Pcy�����2�f���wv@'��YZ\�����t ��!��CU6%���o��7 ��#F˷0�ݎ���Y�=�s�����վ}�)��Cw�S����I��v@ְ�P���s���l�>�kX?7GT�>z��������PZ�R�%��!�Ql�"�}�����O0'�P�� �����K�������koiS�H�/UB*����,��'g=�Y�p��:rOY�ي�/����"�j��`�ɣ��_��A]>�kF��L�7�}�������Z��~㕗�.v�Z�h��	hI����m�Я��0&F�r`�d�Ġ�W��X]=�}�q��5�9%8U�
�@�t�t���IA:�VΈ�)�&u��'�:�F���g.�##Mq$����H��YX����(m�"��LwO"�@�i��1$�B���d�[�`a��1��ȷ#f�n���w�@+ѓ�З���5�������c���5�_kȵW6��J�����nR�6���@T�T+ɀ�3;�T['ǰ}�ǘ���C��P�Ƒc䟷�8������ױ��.ς_:*�K�n�>�e0c|���D�X�Y��o�¶m���X�P�F�*��se�X6\�B#��Q��.�!�A�V{LK�l�Kl��e{}씨f�t0x/������t�xS=:K<�Z�Rmt6pϻʔ�s��������<{�frlFI�#�#�ސ���þ��W�|����p'g�4�����0Y�aU1O Y^Q֙1��ǐ��cG%�? nΑ?&1��E�.H�!�~+J�h��_$��׾��ы�|/M>���_�u��i���,��|ߕ����$�ꈀGev:q�n��n\ӧu�e&����8~�0Z'��-�q�DEӳ�28���X	#,�^EC����2Â�L[�$�ɋ��J�:�֡���kSԹ�Ѻ�����/>Oy��2�GӖW��Ѱ�z�S3v�L�($��Lw9����04Q��v�|��#ÎV�{��ҁ!7Y<rJ�U0��$Z���-��;���'d��>&�O�`>�J���Xq�F�#��չ�J��1e�V�n���_�en#��1��ɴ���s�v]����0^:�f��D6P� ���cU5�[��r��b��\�����v��VgΤ������%x�~���It��er���C��1�ǹ�c��3l�d�;D��>=o�Q�sI� >�,	t�]u���/��^gy@�w
2�>{^֛�}��Z�O��B�0)��˗�s5�e'#H\�ɵ^�38�d�����H��q�������<����a���A�����D�8���ð�^�_�ʒ�����q�vN����u�y�l�?���z�/��P>�$�)u���~��� õ;����m���ր�[��?>x�]����}��lþ7bn�~��y����)�\]��=��:/���8v�mt�ۦ-���{� ��+Kp]��I�4@	� 	Ё�D#�b�T�.3]������������������������j�RI��,E�D�  � �޽|���{�{_&H�U"����Hf"�w�=�ܳ��fm��at�:��x��_�'Tn��c��%`�6�P�?�?�!	o�HXF��MYJ�U3fY�A�Ik3>����7����c�6�ޛ��а��\��1>��f@W�N���X�$�]W�ӺJ�b��$��+C��s&�Nl��9Ĩ���G�-Th�Į
I(�Sf�1<��M�pF��>�X��'����UWr��	o�����ζB���$[[S�a7��%����r��ُ5����賹V�%��i# =�4�U��0���}a�z"��2��9=���r�g���N\�5r�i9��`���ev� b��z�kc���Q�k�C_:��[�41�)Mk':�'�A$`�q2�=���N�>�
]��?�j��!J��t,ϣ)һId�\%=���5�+�g�ں��ݻ�J^^ܳ��>v&��~��BO��"�'�fC,е�qt4��y6x��k��*	�_�X��
����`�6��0����Y��v��{|b��[���ޅg�6;0#��a�nތJ� mX�$�1�3cN���<��Ge3���C{q��%�?g���}�(z'�a��w����f7;��t��ߍ���ӡ%셓lbb�)�$��%�^]eG�b�IN��Xn���a�+�&r��b�R/L��T*��3�0�����9a��Z�����(��C =�U;U�ԥ-9˚��t����F|����c����K�M�Êi| [5K	b�,m������V��6�H6﹆�a��R.I~�/Kɥ'ri��y����0�����j��Μ
��d���n؆�?�m��ŋ�X�p�X+$\
��'�6,>�w��v�c bFIb��$?�<,�2�H4΋d�0�����y�[��H�\�X�jO
X2�E�d��I����@b�m)9�$Nj���p�σ�n�M̜\*-�S1�G� �6Lյ䃴OJ������Ib����z@K�.Q�̰!��B-�z+ɇ����QZ;��'��bvf�ߛ@~�lݹ���p���p/_�[� ����N�7�X󈿼&����+lO,ќ��q��} �b3��X�[|�I���E�"Ԭ0�m���#m��E"�Ck\ZCF��Ӌ:'t������{׈�UK#����aZ��5ب�c����R?���7�K��x��B1���1|��I8n9���yh��Se|�Ҥ4�'N�b�mB���f.5��f�7�(���q*ʢ}�u�ϊ��*�B�����yf�r�,\b��-��I�3�ę|��\B�Dͥ�+3^n�
���^ʣL�=<�6`+�X}Ly1f�����C�F��cg\�iC6|�e.�S�ǘx�}���0�v-n?|?�C�t�$�I�$!���R7���-W��b�3'3%�_-I��q��ă�^A�7�(i����'C2�e�܍�'Pqd��������1d�p��%V��
4�g�#C�̞6���-1i6�8=�}��q��b���6��ڗ�u��{rS���q�\��'��jMiu������%H�t1Jx�X��ׂ�V(Ŀ�z����l����d|�&7��$Nr+�pb�[�`��Y�}���5|�#�7r%X�F1�"z��aG��de��� Zh�W�:ߥ��=��'���Xu���c�o��Â�Gl��$�l=�����ka�Eb�gWk&��F�L&�D�@ư��*��g%�F�ho��5��\��)ת�[(U����)��a6qqvŦ�5���o�M."�"��1q�?�.�V��e��U�3�W2�Jٯ {`H]��d2ii�Q����e��Y�9��T��H]t" B�/��
g7{ZKu�l�����dH���,A�DELD��_K�Y�6]i�A�s�>�#P�'ھ��G�������(2��r��:��f�ڰ��賿��Ͽ�H@����#� Peo���*�=���c�
ſd�f�	�6����I2�#��ZBr�v."����u��>�?�˧�c}6��D�%v�Y:��j��+�*	�D4Z0b��JT�8��vƆ�t��T�I����>K���DgW։��׺Ip��k�\~�_�rO%�M2nD���Ј�����V1�d��9Cl�E�MC�yh��א�P��i=`�jl��E�$�����n.a���q&��=ڇ�=��ݷ�Z-A���ه�3�љ�D��\� ��H5A��q��'�������t��ѳ�z���*�����7����f�9if�ohx�?���~�8u��6m2�@�	�f��"6�D^?�
�c$5־���e7>7G�>T)����]i� �����.˦���Xy.��@��0%�>8ߩ/��s7�M)y`�mK{QM@]�Xv���ѿ%�n*7���0ѹ�>K_9�إ�b�
�uuެN8w��0&u�\6ŭ/97@%����J��1���v^a�I����9V��g!Jz��F����)Ľet��0c�����W�f�@��������;3=;M�i^zbk4�6��g��9��	�X1�C(i�D�%s��v��_��Ο?��>��-[E9I�;��X?Gݸż��a��1x�޺pU�(fU��s<,��J<Z�<��)��L>'��l����LZ�N�T�Ny�\��
g����)=�z�ˉo���H�w>�+����1�˽i����%��{���4ӝ�+�Y�F�&�W��k��X�Z�Wߴ$���oT�v���i�b�X/I�A?�`����'��f���ݍ�3_�N�|)21qnk�Q��n�^����#��$aV�0�P�L}Ʀv�?r��}z�Y6漃Q�,����~������ţ�y��p���XK��r��%�-c�z+�\��y`�N����[��h�{��c
����IM��b��24�,..��h"G�ds�&�`şC[��p��c�]$K���Ҝȃ27j^�-t���7�\�5�5��eP��`(@��k���j�$,�s�p��r��$$��H�ԥyiѼg�y$�|̽��8�-�ݳ|���Hʩ�{�������ʹιT��m> m� B���ሬ(� ��ҤY
�W�VVZ�����/=�I��ќ���A#C-Տ���������*eؙ,7�V3���G������d����K��O~"�F�Ƥ.>"��ݞaQ�Py ؕ�}N���;�D���Q;uB<.�ȆK�<�&gE=_��D�_<қ��.����%I%n���.+6)AS�>�f�NV��H���Z�� �ĝ��u_J�T���1Xsu���x�ܫsO�|���ع6�����8%�����!UN%*��)�|���/��x�"�ω�N!+BI�	�/Oai���_?�Қ�ܗA���=��uf86�:2�*
AL롍�|)3�6���5��v-W�&��[��q���;s��;�ML�~�=75:�U;?��x��t�8$m���&mJ����o#����)\�r[���q!�O�J�3���0L�������'�K�I�r#���L���(�������<��ب�K�Qz�8���F��PEIV�<b.�# P���[cj+���#B���D[��bSLQ��;�\��C�>�%�3T{Uf��U�I���M؛���A��2 eW����Zj�|.G�c��͋���%.-�u��J=b�Y���Ae�&�ȅ����ft��$.��,f�1��;��O��#�m�Z-����,�-��;Gq��_�;}�ƍۀl��,Tپ~�h�+�G��\���6�mFoO?Ҷx:�nǇX⑈�Hܘ�F�ץ^��Ǧ����铨�0�����j���H�2��}�A�՜\�'�����
l��F���A�׬�,��)�G*�_K�W��k*G�Bq��,Ԓd/E��LƑ��}`� ���a#�����á*14��&!�P�֗-V�7�c�e�0M����e����4�AH_�t�x��4*J��1&	}jW�p�;��Z�#k�c��+@����~���g.B�]�9�����ȸ�f��H�m<R���� ���|O9!s��ߚc�o�����[� �
¬�h�i@ҜB�i�%��q��r�b��	��mT�E)�ŕs�b��Dl��6��6A��M�;��lm��?�zc(�	Ȍ��^n��M��wi#�#�H��'[}wo��-�^��6���������ؙ�
k��ϊcv6�\�!2����Y�Va�kJ3�er�a�k(�s"�*_�
���oX����E�xY�&-J�N(�^���x���"<��ub�Y)e���e�]aM�d���R�K����3ffl&{�*8ҒVqݳ�������Ǝ<	md#<�w��`�Xo�ܧ\ �P�^͌�#+�je��v��%��Z����?�!l��b�m:N�P��/`p�V���{�f�����#cq���b�mwa��-"t�����\]5	1-]��I��ݸ:mGq��0wކ�K�:*l��%�_4繫���к��������bZ�b!�7�]񬝟����L�P��슖�=uKa���sT0��^���ܙ�� �7��PIx�dǆ�xQ87�Y<��bu�hj�8(V�x
�7�r��W�Z����/���_-i[ik�1�U�Y�M�{�y�5v�
%��K/o�Okyz~#_ލ������h��o���Kk=�oK2�"�=�/]�P!g_��i�!ү�u�d$etf髱�[q��-8N<󄰀&�*�����y��zugM��H誻׀[�@3��+�n�o���{�b��1��a�Y��`
(U�12�V��ZӳX��pw�槮��р��bmn'ڢcu��j�E�������"�=�%�މ_|�?�ʥ8^��p��*�d�nEn��	]�.X�YƲ�8dld���byd6�u�\�m�M^���nUF�򧏧6�-KS@����c��'�M2"8���:t��7�(��'mUca�U�g&V��ɩ�|?ڄ� �i�R����g+)VS)�r�N�њMېݴz�B��KD�!Jf*'Lu�ҹ<w�2y�ˉT�0��g8��Vï�]����[	�������t��i�S�}��;���S0vn����ڼ�>����MX��o�w���ufg\#��kՓN;)�s��r�b��
�����f0Bȗ�M�l�87'��NVj�C�������IV�c ���2�����[rWS	����ە�1��Cb�d�zQ�0��A�؎|>/F��H�f�P'`N�̪hR��Y�r���k���`e�����ӰA�c�KW]K�Q�ŧ���;!}֓�!���f���W��&$p,%ސ�a_��,�u�.��t^=��F�R^J�Ȧm��L���2 -�5�ήk��E�ű~!
��T�U��[q��-8z�{T�T����u��v�0�����!f�m\��W.��/�Ǧ?�*��E,^�*���͂D�#���*Ī2�Y�DG�OC��KĚ�L�����%��	NĤ��ӗ1e1\@ax����[L��6����u�Zt�R΂��"v]U��	d�X8�v.�PΘ����-.O������3[�%��Y��S<QӤ�Tw����(���&��x|�t}�1�c �cvZ-2nh�t����G�J�bJk���M��bu�@WR�� >���\���C����諲��ʧ,=ID[N�	�ʤnA�+��C�ť�^�����z5ҹf�(��is��ļ�Ϝx��8���1t��(�����Iچr4p\VSB9�8i��.��/���	*;wbh�.\�:�������4�{�̜���h�k���3���.�����iH��j+�u�NN#@�g�i\��J}.Vb:�x��p6}@s"�k����-�qx~-i�B���|CK�5?dt;�a9��^�Gl��\��y���tMW�P��_`�G�c�� ���l d0��B�1�lz5��r���� ��/�s����ރ}f����l����8��=��W^��u�*��b��7����ns-�fE��Y�{�jgKv%�AC��V��fa�)p��`�m�~�0��k;��̄ݹKKuL�����Č�1	?	���1y��x#`u2�)ܔ�ؔ7>�j�G~�����ǯa��{����>p;���ŗ_���s6�s�6\:ױ��)�f���A�F��﹜�R[^"�I d���^@�ωhC�\)�	
�$�߼�l��d�Kc�"�D�M� ��.���wfjZ��4?��3�"'����m�T&uĹF,,��Xs��v&�	:�M_z ��[��a�Ϛ��r��X������+�##Jz�$=`|��/��W��@ij
C��^:A��4_�/�@�[~ڢ#��k˲���@�w0yu
s5������e^,��s�W�
L����/O �L���������̟:��'Oa�ޓ����sg���R~�C��/�9dC�c�&���u}ӡi�vY�g U4�Mߕ�7v��3s�/�3�\�Aǯ���Ul�������\9ّ�����]���C��'���T/��H�R���r���OG�R��Ҡ�"����"ȶ����(m�@�������;t���B�>��|��^�Vk�aݷ�_������s
m��D�j,����~��xew �>{)��2�ZۆLSs�e�� )�axw����9nا��=��K�������o����fji���U��cU-:���>Y鼩q���:1���5��M�fb��qT�a�K�!x����by���c��0�ȣ(lڌ��_C��7�_�@��.�X��w�(�}bM:fܦ��e�\F�QG��L$A�5����̬0�Wd�ƪ�ȧL}Wn͛�Az��&�͜��1d?�U�PC�2m�u�ɜ1 q΂����iǵ$ю��	��F�@�[�Vv�@���:	���RğH�%��4�)J���b&k�V����w�_d�m�fPl����t���%�qz��)�և۔�hE��L�����qL����m�=�$́~�d$ľM�`++LX�*[ɖc	�����:�
c�0z�!�y�
fi=n-��U�N��6�����
�Y�]��Fb�Ix�{�VvN��1��I��E�m)� �n�2��.1_�b�~R�KI"�e��U8$Rɜi�C��3&�*d�'X����*J�%��Jk����kik�
���hJ��/�r�^h�6 E6Di��5�9撇�ցV�Ўjj4_�9t����kn�@�ԏ�<^"S�m�ϐ��k�X��X�[h\#vήK��8~l�a�s��yb�v���K,/�o���b�V���t!���<Y֓?{����ލ1�v���<��[(K"�jY��viot:R�l������-Y[ubT��&��,��W i��q_޶秦q��"����c(m�Ła,mڈ��_�̹���s���ؽ�/Įx *�Ė-J�g�7�-ٴ,��8C���iݎ�������b�n-�gZ1�~^��2p,-T1p��(i��+��c��f�0�d�g�Uu�F�?��͹�:�������\������;m(/'�Kw0�*s[t����,��ז�>��D���Bb�n�z�tf��}�%B����;��b���t�<�8�BE��!e�1���	L�]�s-�D�q�Ar��12��f0��0�d�ж��y�A �Ii��jҽ�TI`������̍e���jJ�WV�^��Z����\[ @�X�Ԑ���;h����b-�Std��Ԛ���)A�D@G�p3�+3߻�U���R����x�Z���sAsoeT�W�q�Ա�g�y�����Ǳ������5�	���^�����g�m�+K��Z	�Ș:�&BˏEa���3V��=���3s����8�q�+���6��%.s��Ze��RN�2h�&sz����7� �g������[�~�������,��yz�[m�>��z��&@opͱ�Ԑ�`q	��	ؓ�	t)w��z˦����}����W}
�m�ѻg�|�;�@v+��y\���b��9DKJE7"��9M���f�h�
y8�!��MciiIp|ߐ�Z"ՙjr���?c��I����d/VRa��%�*IW.�b��mV��s�)"-�F�r�Z��c�
_�$#+������,|npC�1Ol������_��b) ��lPu��Ɗ�r��o�ٟ�8��>{}�*����]$
��}	�$�ò�^ʴCјgW�ej[���`�Z|�!�#������ݷq�Xb��J�,i����ĸ9�,��!3��|�.��0)Z
b�����Z��wc�b !�����Z��I��H��^��;��AB �%%r���d�r�f����-����ђ>�z�Vvs$���7���܉8���u����;K֬ʈؿ�e�z�N���dd�:�.3��N��ͣ���K�$;��w��g��4����|����hꏛq|5��8up�k���*c�o�Q�D8��Yh��̉C���x�0�m�,,
"qU���Lw9���2`�9��q���َD��&P���sW0�gzw�D?���F�2��[j��g���6�&f�\�a��E�KبQ�Ĩw\��`t��|���J	��Թ̍v��ڝ1���{�cpg��{�NC���G�J���7�(��'^0��ev�s�n�tJ �U�ߺ�(v}tD+z���hO�>�'�1k�9���x�%�J�;�ܵ�6$��:n�I,���i��ELF�Os�@Vgd[����#�X6ש[�ȯ��������GWLT��%�k�$��&�]�oڊ�w݋�|�w�j,�q�K�8k��T�i~Cv��ӜF}y��n�� e�i���gF�����ǡ���Ӝ��|��KZ���L��1$�ݻ2����e�;p �.�����?b��eH�z���_���(��)�[��ڵD�i;]	}@�s�	�Ga����
��p����b��]a)ל����s�zC��3ܪ��#K�D!�W@'R��=R��T���.V��k�f���X��!K,Ҷ�R�4�_�J���I��(QQ4�	�7��1�Ⱥ�O^H@�=��8�[�r�O0Y�!�͈��ҳȘ���E3bi���\���^C���{������Nk3d�'�1}�XM����*��㽧�,�pܸ#�}M�bO�m�Z���P�d�.�[�ڌ�E4#z=A9G �enLb�B}v��%z�-O5)�����q��{M/
#�(UKR*�P[R�2��Itf� ��衶[�ú��"����N���9~"^A���w݉፣��~o?�_�n� ������O��_��?�	�����P#�?@��p�B�I"Z��$��b�U�^őuY�z�b��o�u�a|*����W�Q���ԝ�MeJ���v�����v�ď,,e3�� ��aB��	j�ʥpv9���fBe�K�%4Mbº��%	s�w�e^ۘ�to��605���
�����L��e]wbd�)��җ2&�4jhq]�
�@ў�P,�C;�~�K�lC�u����ڒ��]߿�L+P���s΁��*+���{�����&/.a�ڇz��j��2���� �J+�o��d��8��
���4��E����)F����sR�����Ic�E�y0ETF5v��4��;���X)2��t~ơ��b��Z=����煈@�9�ܳ���ՄǤ{.U�~Zk�о14��{�@Ϧ��O\�ɗ^@Q�lvZ��Gĳ��-{\�{�����ay_2h5�X_�X�[`T-���=�N�km���\��.,Ifz�v�"�Ӧ����l��]��f�bL�['�\7����˵�?9N~������Zp�j���0������dq&t�\��w��M�X���1VƯ^x�����I��c���)���}�`�й:��sP^��]��cWgQ��mx�0��mÃ۶b��wq�;�Õ�^E@细�˒�6_1/h���"g��$�\D=&�z��Xo��?J&����T�l9��\N�� ��gH�S�Nv��%bC��z	 5P����ULa�L��?]W���b��fC��?�̌���X/7U��Ͷ[8N�E�Y6����;{\D�/�<��u|��w����w���#Fn��in5xĦO����3�����b%�ۖ�Lع"�rͦ�J�l��g�g�7<�w._BW4pkπ��u���F��GS%��5��n�n<99��s+�ً��+7�&�Xҕsb)Os���$��g�[��'7�1�K�TIo�c�����0���Г�)���;��8ʘ�r��X�/Pu��M��ˀ��6�G��_�����F���{Q��0���B����p���Gg|dqf�2E���\�{�0��\Ҥ�)�Z�~�a���K�"�*��CDdh�!֡�a0���C�-:d�&����X��WAuh����Q)@#0\`7/m��R����:����7cI�ѹ�1��K!fWd(%<-��5�F��&~��6Y�>m&�����ϵ�0>�;��O1�m;���X�O��ƾ�$���������ĥ�8��}0�X�v�=�3��q�_>������=�������.�/�0H�i�� ̗(�F� �P	�Tr�.�~�$��ˣR,On�?h����'���7���MU����X�C4+���c�I?z����$	.�|�Q+1"��&~���j�А+b���x���kX_����)���M���������
m�kGF���صy-�����ԏ~��'0f��Y� ^|�W�m��p�$ ���5D�<@U�g��?#:�����q��W15SCo���ΐW�,��/��:l˓�+����,�(V��>�Xx���K-C@ђ�h1�B�f�/�rP	�<����� އ��n�*n�A�����D�6dA��Ü�ɼ�)\H	)�y��bŧ%�ņjT�Z2}�x �������߭�
2;���ً���X���F!�\��{aa�pZ �qq`�M�h���(��B��cc>i-rU���6V�M�*����xR����B�sG���d8�u8��f�&��Ă��<2$��w�f�V�gQ�6�����h�O�>>���"�"1y���hӆ��ݝ���&ĐK��=)v=w�]n�����Flܾv�J�r��o�WTG�L���K�U�Un۾�6���gp��W<�`\i���Ʊ�8IV�A|>l��0��ƶ`h�m����X�tW�5�袊�Scяmh�m�V�I���q�!��|��1nl4��j�k��k����7�k�K��][P�s?�o.�eAu��C�&���媼��5�˹�i����kr^�d�+�6�X"�Z\3�=��	Jlu�F�ȑ˖�y���l.W��F��#��tδ��t���Qo��z=�����T�oG��p#�����\M���%y��3���7m��ę�u��A��go� ��r><����$:�a(�fܫ������f&��Ri��E��K����<���-��v����X���P�Z��+u<�G������;������B��%��}�$�5�;��l=�FH���,�� �/:\��i#9��a���dP�<��'O�46��};1t�=_|���Y�7F��A����+���ժ�����U2��f�HF��C�b�j]�6V�ǿ���,��}.s����(���浛����k;��A`�D��/.ڈ}D�8g7�wk����"36���N��µI��Ț����4�j�����'zҞ��H?l:���Gg��g���Ff�������5��ѱ������p��F�1hC��Nb���[o�9ep��\����>��'��| f�(
p�ȍ7��N	۾�.]�䛯���4f�.����o��p��$���������K�Y)�"��o���i
���Hۦ-u�K\O?2@,�0��5���FV�cc�����Nc�� y$���v��B	����
���E�T��[ݶY���m��k�~vEs�Q��>K[!J�롭3��m����dH� �W�z�	,^�����B�^�u웳%�!�p��7��'�V��R�Cj�99/QYC�����q�,��.Yl�s}�;�8'�>�@Wez�+��
�n+B<G����y�.�
̥���po�FK2��/�lC�K���6�\f(�I���q�#���kAE�R��u��BUKJ���y]$����^�Eω��?/�x���J�&�{L��Qޣ���/�z�A?���`�G�B�%�09u�p Y��:���Pr$4Aϯ�i����b���-���O��/r.�G��c�J�~�cп�Q�-Ur�4t���G���]��}FL�l2��$v��Ͼo ���U4�6�2�:=�-7�mrgbW%��dYF�Bi�:�f��k/O��o��؂�襍���A�]�"�WJt�}#��Z����6�k�~o^����ޏ�Aa�l��o���[׋ ˹7���;G�{lz�����i�����(�
�R� �>���8�܋��v��ğ�K�߶��`��ط��s�� 4��,L;7v���c���)��?$�c5:C��Ln�&4���,3�M5N��j	[C�T�Բi&���Pb>&Rb�I�8-q�s�"ojR�n�����[���{'�B.��q�PK�a�\��`��Q�o�o019�K�/�|��S'$g�{WGdPqI���ҽ��9?�E�.d��|Q>�[�Ip�v�r���0�k1�� ��R�8��s���Q���k/��}=ʥ��W�N���;���gC���7}Z��	������ޓ]���ƵksX��#�J �F�0�.�_S�R�����N�W�;V��P���Ӝ/�C�ݢ瀵���;����P��~&ni:͕ٕ��$���*��}��4�R����ݴ�4�#=Qu�D���0X�݂�kqW���c��F� K^��d�K�kӹx	�s��Ե�h�:�}�k�ٵG��%�
�C�k_����$�?�)�^��	�����p�豊���*���y���N�zd�.������_{���\eH[e����8�W!ky�����"v?�(�m�X���ݭ�ZMg'WE�ҏB�����j�����ػC �[�@a
Ch^�F��5:�O�nCoF��T��b����T"Z���������`mn�~��X��(z݁�#b��M,?���)�y�8��I��e�@���/=���K���ʈkuL�~g�"��-2&l'�z����p�_��=1�������� �'ϐ���(33�؉��{l�BxI&��{OD�H��#EYX��+�	pC6ʕnv��N�]I����,����fʐM@â2'��<'�q���d|V۳��#���}�v��@�*���@���=%t���ŭ�®U������t]k7m@eM�%�Xr'������4i
��(34���c��1�Lg��\?�$�	D������o�3��
�p���8��"��1�2���۠��K�|����h��t%�^"s+&��-!�*�Đm�K�Nci~e��{X������"�6���Ī9��l���|�)�3��K6�E�EO�|k�7�I�X42@��â16�g��uǪ�]W.l���$i��J�[9҄ț�Otǋ��w��ȫ�H��X�o������XA�k۱U. K1�*�����}�Z��e�%J6�c�׿F��i\WĆH��uk��M,�<�K��1��4˖gB�i�<�w�s[��C�~�
���*}Z�-#@�Z�x���*�A�YM��X��Vtދ��B��7@O�G���f��C��ۅ�zKܶ��a�X����n݃B��6=���6�Y�k����V�.	T9����(�
�1i�����,4�8ޛd%1p��F����"�Թ��۱Z\=q
'�;���'�����r�^�9��n\�\�h�����{g��G����z5�x�y�|p��ĺ��пq�_~�=�3����(�b螻P��v\7�ډ��=�"��1�Ǝ���Sj�[���mvGj3M .�"�
�ca��D�L��)uk��l�R9I�ZU��G�i�m4��0�XW,�9R�͊��DXR�բ7O�ܮݺ�ƍ 1u��궃�C�!.PKg�wΓP.xq,'�k�z�������D�s#�Ұ#�m���a�oK �<>~^7���9:ǜ���f�ߖ\��� �3g0H�W��@�mS�d8]�9�X�E����0��N/U0�w7N�8�6���n|���F�7�xءg���"���Ȓ���-vs(
"Ӧ{���*	�R�us��9��q������ 2@Ϳ�?���߿?|��_���
yv6`OK�ď~Њ4���!e����e��/���3jﾍΙ�0�G1O/�>9)�vlވ��i�W�cK/���2�
&�ڇ4+{��}iذk��z����ګ��wï����{��0�?�~���B���}��4}�45f6==������kX�4���ص�m�+S��(�蒤�L�=CC��s�15��G�EF�ɗɠ4���,���07>-�t+���p���Չ�g#�m˧]�c�1��X�6��L5�;}����K�|�[���ۋ��1{�:N?w3��/?�!�wbl9�[\�3���Y�;���!b�����7B쳉��^��^y. �:���1�'O���c��E8Z9�6\2t2pI֥	E�6� N�i�׊0��}�J�b�y��ݗh"�B�O���|,�t��h�s�0�����s�� u��+��o�t�&êz��}�a`h@e���]5yCM�ʓ��]Tm�8r�t�E�JX.������!���Õ�[]���IZI����yX��k�|['������@\��:71�KG�����K����L=FI .��(J��̲��<�!J�VF>���}젵iw:Ȱ[(t̹E�OF� �PH{��d��:��Kܜ�굥%���,���H��B�����\Db��e-��S��[x���^��Qy lpsnI&�����I�dO͏�v��B^�k���|,�F�{oۉ
���8�N#��@��Mƽ3������Үz�X3~���G�n�q��E痥g�C�`��au|~c�?��֓�#�%mbf�w|�k����;avnm݁�M���A��@�ڋM�a`�zbx���ψ{��8���*�����&֨�Ѓ���|��%���T���C8��8�����& 4ԅ����g�c3AS��Z���+��,�2m2W�<�����{�~����X�-4��ib�צhSX#n;�\��v�����N�Z��<�$�'�Jkr_9�cϽ���oは=���{��c�N�ŵ�����Oh8Z(�j��s��1��8U�ԗ��.;[���e�����k����G�@������xsIu@Z���w�#@
Tg+n[9����pvmr�Δ�d;6�3��f���ּ�o�宩������g�4G��@��]�O����D:X�K5��=�H���� n��v�,�d�M�;�`~f�$�q��t�bV�&��$ƝV0�r\=n�Ъey�Oc���ܝ�^�[�;�=骧%��*�@̵��K6���VG��h{-����	}�h�����8ɢ�����9��3"�Þ�H��B����!�]Q"��$l�d4���Z���]2��|�m`��=��?�YD����г76�c�Wў�N�A���箐��
0�)䦃�CESN���pe!wK��>��Ux����Σh��pvx�[ݻB��jVq��Z���hs*m�m���=�l��b���ȕhC�͍c�i����F /j��"�B�3S�X�Mq#���&`߾a}�7b�W�i3�nL�6T%7qY+H1�Xo�}����h�}��+b]���*N�?�3�m\��۸�kOc�=wc�]�q�ݺR��	h��$��x��m܌u�ѦP�����f�&�RO��ױ{t^�����_ᾯ>��}���c'6�����k��\:�����:�-h��u��8��@�Je�(UFOkٵDYT�N�BN8t��OW��zt��
d,��_�x(����ˋulz�Q�=|�[��7�3�YO��b�X�<�]��ղDU\�t���[�dl��:t�i���rőRM�9��'5��)�᳷���eC���dT�M�`��8�6�JI�/bQ��Y;5�)���ǂh��\a�6`�A���������o{p��ڢ�mjV�|=�J3�[�#�Y�ǟ�*qn iI�����6�#��bDIԕz�+X��>����*�=����Phh�'���rN=�U�*?�P��s�i�r�K��w������Wq��5���!T�P�m;꿸�R=&ÿNK�F��j��L{K=���B;A�|ɧ��"�����ױ:>��
����+`�� Ԍ0���1ڦ7�!b�#�� �n�&Td&B�.4�`v��v��s6t�1:�M��nr-�T73����C,Vұhs�k�q��W����]��%�R���%Q\��2��!�tb�ČvlY�:}fPk��܇�5�
f�N��_�Z���3_A�@;ȱ�5�ћǶ�v�����?���	�װ�����*����4��>�}.bi�:^��g��w�۹	���6���Y��q��?ƕ��� �Y���� �>��܍4�7�@S]U�i���J)~�e`A#b�1?��%RyK��7V����;��XJ3�%��C����� zj'*s��Z�\t۱"���K֗m�B�ۗ�-P�uY������Z�;f�q"'�����	@�Pi���:��������ΜU�Y[<
Q��`�kd �д$C�V�CkY�H"\v�V��ۃ���EI��l�������e�P��qK� ��2h8n����1�y���\��'Y��M�t�d��#���p�0v)�>�yXi,'�9��Wk�2U��������1r�[f��'f1~qA�7���}/�g>������^2��y��͒����;�Ѵ{驛�Cv8�Ƥ�-�V��7V�sǞ��X��Υ�Ѓhׂ��L�6(�%��Ӷ�ͫ�*�X���㻰�9��Y� �nF �Cφ�Ř.������$mP�E%o�J3X;��J��I�O�X�Jƴ']I8���nh�Їn!�Y0e# ��6QW����ן>���w0��i>t�M��h���C�}����1���~���������(l&K�J�%��lLO��S�0|��� �]���^y�M�e�(r�wb�ڃI���_���\�������pm�SB��X���۝&��M��6ͭ�v|.�"h���NUt�4@��qhnf�R,b�EϾ��ʍ��Ҥ���
�~��\u�X�����Z���j�+w���8J|�?�tn���t�Y/+C3���䶣��%���w��lC�ĺ�	�ʛa���S8!1�5�ٺH�sI���PmW �C����R'?��x��5���"�	H8|�(��rfz&W"�x��C��>?�[ka.�jZ�]���%B�l� qKG��^�ҵe���qsa���8��M������v�ʼJ�&C��JI�S
��w��;��<Wf�u�?J\�0vS�H5YӭFޕ�����<|6�ա>�{k��c��>=Nsm�oӞRȀ}hmX��մ���Ny���N��h�B��9Vg�s/?y�KJ�&8�/#��dd?M���R�Ӭ ��&f�!�`��k�k4Ѫ/Sj���&������`W.Y�J�n9o�{����DR7�<%`�nZ��5�6W��[LN%341_�D1�Ks.<6�=Rs��L'o�,�17'�H&KP6�!Іn���&�FU������<y�;���wa��#�m���y�}\y�*���ڒ�2�ͭ:�V現�F��?�&n{�l�����֮e*��ׯ���O���ԫ�c�\s+q�j7edڍ�l�X��˝7RM�q3�C���O��	A����ĭv����֢��0
�����ǎ����a�6��]֨�<�GNS�����	S�b�Z�a�P-J�(I������Mq+�SK��S��H�Rn�B�I�]���U�^o��~��e�F�5�9�`�Ѡ����7�J]8Wr؁5�"OX���)���DqȮ]1����N�|E�JEht��L�I6~&��EPf`hX1vN��T��/�zf�Q(ƃ+N<i��/<\j�����g<V6fI����=VMe�D��=F�*@���>z$N�eK��%01
����G����1�d��fq��_�⯏�B$�B7��X@5_E_���B��a����l�=H�r���K2~����֗W3�?��
��(��+��0LV��9ď���N���C�p�l�fNׯ!��B��E��+�1W%�+�#�����W��3U���h���:�y� <�{αc�X-��iS0dcm�S��1X�:4�z�E�6�^.Gb�3b�m�3�m��k�,��H�%@����F"��4Fhm��t�BC��{1s}��l}�J��Ŗ��fߐ:9]w��p��	���n��ɓ�x�4~�Ily�>h�,���ۄ��Z���YĞ�(oC��Ø>�>:�s��~�[}�?�	��d�����(T�r�+�d78�
�>Y���&}�2�r6ÑNf�Z��}Ã�am݄0_��2�5o��q$���Uz?O�V����k�$]	IK�]~��J���H�a��X5-��Z�M���9�[���!]���z�5p��(��@�|/;֔_�_�L�RoV�(ތȋ%�CO��r=x�q"�U���#����p�Wo�z��g�04%́����y���LFU	d�(�+h�������܈Ų��O�s�K�<��>^�ЗY=��E���1��P��f��M� ���h�m�\̝��3�E�9�^2ʳd��:�e�+d�M]��l�����}sz�M��h���h-u��dh/x��{p��Ռ��z���0^ v��2��4'��Y����jYbHY����b�6�5��E���X���v-���q,\#���	q,q�[��=�1�6� Щ/"\�Qs�~���+V?m���eg�Xj��$ ���
�p��j��A,����Yo�yq	�^�/���F�)�i��� F_*�Ld�JC��'���ŷ��篿��}8�g��{"���ju����/����3���o�g	ܙ�<�8�\��|��;��s�4_{6c�xQ��[���~��{^��7�
�u���I��7����U f.�)�	���f������A��"����>t'�lF��&�L=�)_�M�'[�0p-y���@OS����t6C���Z>w��w��aq���^)�KB�#{q��E[C�h�b�z�n�n�4���Br:g�'Jy.�;�7�'��G��W�~��
	�4`Hٙ�	�R�ϱ{s�:�|�1�ûo��Z���V��0oՇ�'p7��Ɋ��Sy� ������=�A�u�4h+�n��`��I^�����b$�[nn���wc�+'�KS��q�{̿�2�SK�kĘ�i`����]{qϿ�]%��Q~�v}�Zh�J��x��da�;s�֕+a�ƶ
5��X���a0;g�M�l�F�����u�}xMl9V+��:m`�f%�"=gK׮��5mt������V��#@��{4D/�g`�RYb�K�3h,��
0;5.�N�A�u��'b,6,TJ��3s58�2��O0u�*����������,�>�յ;mb���2�9b�����Ѓ�	s������ڡ#ر)q?N��ˁ�p��@}]]Ǖ�'���X�M��g'
���9=���Y\x�-�8{{y9���M�V�s�"��mnf�M:3#.k��1�rG��-����@��/ga��
YN�Q�k'.x�A�-��B=1��:
�*��*��d��k������'�p����\��$3U���&	�G�Q���Д�\K��V���q��ɧtĉ�7�9�L�Ԃ�ݨہ��:�/9��ܛ�h΃�kI'82z�K?N\���+��`u�47O6�'�S�q(b3��`Á�3�q�9��B���?u��X:�z�L7+	Uk#4�@�FFВ?Z��e9�e��G�<���o��#Nؔ�}���xe��oZ�S��}�p嫴Y�l<��8杯���ڛ(�%�
Fw�Bf�>��,�=���KW0}�,�N ��J{�"�tܲnT����G�󑦟ei�Nȥn~}��8���X��X��x��ԣ�SĠ� ֈQ�5��A-t�����s��c�|3"v]��z��K���g�����ub��.��&K�v�,1՜�wu:-�ĪLn��i"v���@J�8��;QY��N����-{dvk�=�2۷c��Q\��Oў�D�6ʪa������$���},�M��d�Ov���,"r��4��$J�#m�̬i(�!v�g\>uf&�ݲ	�z�Kkp�X��m�0x�.l��Ŗ�P礮[嶦��d1�eo1m>����=_2�%I,!j||�j��>!�q"s�-ץ�S''qя�{�kR������-���S�����>t/���d�E�9l�l�/���O�[w.��v~e�U��ڊ� ˘$�u�b�d,jV�=���?�/������h�����K��a��Fq�vѶ#�������V����>I�괚��Y2���g��ܱׄ�"��f�E�������N��&S��(���ߏ"k���snG�^c�=J|=��	d+ۂ�7^��^�/z,'ߥ1s]�X��؉��$E�qq�ӓ�Dw-u��-Ge�0�!����菞7a�ڎ���A�}@���"����N�a��e����	��m��-�)������_��<i#�s�ڸ�����͎��eFq&
��<��mN.봕��%Z��"m��0���z�fƧp�;?��?�z�����],��h�&ז���0.��p����\̠6?/�V�jN��Ɖy�Z������Ϗ������=���a������3�m���_�9N��gX�����R����g���V3�#I3�n�!#�$g򱜼�{s�OɄ�Rb{����z�6��N���x��d��O=�u�0x�N��EF��Q���cW6m
��R��T !�i��hLMK����d��%�L���2����I�eV�㧃��\"D�������-�N�d�S��n-�����{t�O CHe�J�T��k+9$ANO�X��X��섬�Bv	������W���Kٍ��GI�q�H0��r��֑�Xd�(�.
=����u��,�;M��B�M��H���ƍ�����<ֻa��%g�]��X�,$��<̬M�+R�k@el��sk�d�,��ɞY�*Pb3�������.ޅHT��/�ѵ�t�����<Z�щ������HK��n�d�uC�&yI���t.b��;��4ڇ	�A�܀(�D�'̑!_��ܱ���Ҿq�/``�Cc���fiO��N��(����Ekv��(��;�cŌ�j�'9%��n|�w=� �������ϖ]י�w����~�#�Fι��H�b�(J#[�gl���]�r�?��?��j�l˞��G�HQ�  �  2�ntN/��O�������: �ƚz��^�w߹����V��O�>~7c���g,S�M�殗e��8�Ù�y�$�FQ�hQ�f���S֡�0��dP����1�o���W#���\+���,��J��~2�.U� C[,���.�r�R���W�hu��|��?{�]�N��zN�c���x�Ē�b7|�	L���E�[�ҿ�N�s�\����'���Iz dΑ��b��u%W>��x�Y�rs%u�g*|+Q�-_3�ȏ{�Pw��m$+�H�KX, ��vTo��D������23i" �b�Wr���y��X�K�y	˯��f�c	b�!2j{X�3 PY��;�� &Y�|��l�Z��Ҳ����R,��Q�"�\�徽��"Ny�y�D��GO�5����e����� $����k�A&πა%~�<������Q��Wa���!�3��cʰ���Na�+]�o���wGc�E,�1�kX�r�
���{Ҏ|v������%v��D�<B_ ~Q�¦X�/����i'y�ж�k413ϻ�Yk\AԸ�Uڰ������2�`rw}�Kx��9��{e��d�=��;(�,D[���-�&�y���Y��;7s�I~Ś�/��p�/��q.l�G�
s��o@^|��)�^��;�K�%��Mt,�]�*��z�P�����>~��Щ���J*
z�v\�M�aUd���M�磁'N��?~-Q��bT�Z�_D�")[�e_SB7��0\���r�ň���9���Tɕ>���hc��ç4�9�4k I8ށMd�N�m�w0]����Kx@������[X:s���(�ru�'tԊ�v��@ٽH�Z�^�p����

�P��������2Ѯ��/����[�sk8��K"3S����G�k��/c�U��ݧ��o~�}�x��Xa!�
��ggD(�t���c��ə�đ���]�kZ{�bm�_����m���.Uw�*��@�C\x��~�Ŀ�v=� ��,���/�V�H@16��A>a�� �X�ɩSh	�{��h�x�l:C����q3�[,7�x����}YKyf���@��d��V�᰺ �����Lg�w?�(��m�ٗ�e6
b��2_SfF+5�E)P.n� ��W�o|����Yj�Mb��2On�T��u5��˕tƔ5Ţ<�|ĸԍEV|Y����;>�F5Q�z�簥1���a$J��5��e�T��$.��8"��wE��*j��(�r=*#,�+�	V
�q��q�6g_�|GZfH/��;���[����)f\Vc$��W���~G c`��y6$���	�h�������F�Ohg����=pQ,?�?\�ch��|�O���>2_�}4�AP;�iM9�y���W��G��5��y��/�_��NP��\�J�oQ���(ޕ*��0QmN-g���\���1q,�9���g���~c�G�/=�J�%���W���+M�If f�T����Ja�q��7-}��X|�(�-4�mD}vB�@�T�>K{�@��X�l*�1�K�n�T7u��2�ssX>t��.&ªX9J�*����PݴǞ}	o>�N��j�^��t�{��u�c���p�7���<���y4K.&5��-���.�5S�uJJ�ɑ���H�*	Z:�&UE҄ݶ�V�S�Y�ܹ�gq��q���p�C�`�����k��kO�P��ni'O���������A�1?7܅�4�+�?.�,�h-5y��T�[��h	@�d-ٜf@:X��Y�trF�v;ʛf��z�Yw�v���y�ཪ��-,�4�K�N����������fҋ>�=��NK�8�.�vnI�բ`�F����u'�y���e���-:/��X�L�3�{�|��`��DI��B�ij���3�˼�+�_�C�����N6���}�n�q��9�[�h��B��(E7>�8ƹ���@�t�#�.ʟ�R������D�i"D���Lj�OfX@���ѫ�'TJƇ�#�q&&�N$
���(��_���W��j�GT���u��)���>�y8q
��9F��R��"��;7ȯN|��<�^�=G~6�	�u��]�������t���dN�O�/,u�[�F��&(�\���R2��)
�w��n�̛������ܻ��|���q�T�
��{|w���$��3��]%��>��;H^?��%ƾkrnC,tzD�~^c�[��p�<�b-�J�*��E&'�u��[0}�.�]�W��i}�`�Ă�D�&�e1Ժp�J'SX[@!e�8�0��	�C#�!�	8���,�A*�jG,�>jN��O���yo>��?y7�+h�w���(V�X���p�7/���;(]� ��D��Y]QƱ�g�Z�|d��Y�JH���l�yf���5�m�ҁR��kR�l��`���a�7+_;�S*�����*Ǿ���/����|��OOy��k�N����k�����,�9��X���1�5��3�TFmv#j۷��0�k�kVxI3��F�Uk�B���Ɠ��Rجs
��ªXV�� {���M�����������J?�������Q����~hb�C�:�]�v�8>5]�2�c��c�#��ȿ�&VeO4a�5�B���r��X�,Qc�H$�X����ٵ�g�*cT�n�#��ٱ�|H[���z�ځ
���kn	=����w1 ��۰�GQڱM�}U�sz����w8���vc��X9��F�^m�x��%�K��9��I������[��X�����WW���������^���j�6�i�OS5��R�A���j��E����;r��P�"��8��W1�4�[�LVŒbC9�bz�X�d����0�G���A�5��,Lm�jO��<��b�������n©��4��ݶ]���b���N�n��h%L�{7���B홟���s��U���f�"t�-�@g�4��Ar���P��� `��Trs��� (�ܣ�ń��*�yg��[8��3T��j���((���u��*T�ǋ�@�>�"��@~��\�;K����s�C��i��4��
���艂RE��u�;��s�����}%�q�D�PM�Q�!Nu��[�N�r��Ӣ���*�������9y�����s�О[P�-�fma�W���U����0y�~x;w"kDzϬ�%k�����en+ꎵ�z晉�kIs��5@��f8��{�tO��4���zT�g�Y��/���>*�\�!�*0diˬ�8�~�aJ}n�fY�Ɛ���%Mn����a��p�_h(bҏ����ŭ,F { e�\�$�3{��ro�	g��"�s��o(F���>�0ّvˣ^��*���ív�v+���#�P��S�{���t��Z:����r��g'����JVr������}���W�k)��y[�x�݌u@���w�xH��,1T�b�L�i��(s��"�KI��ͮ��^g��NM�+{d����2o��ȵ���S���DY9P6�ĺ<�h���5�#�HmѼ�Ĳ$�̫/��[�7]uN�s/<�+8�|� ������b%��&�E����ӿ�.�n݂��U\�{_Ǟ;�س���s�@}����)D�.��>=֢�T��Qɴ&�3�����nܓ�I��(Qׅ%J�b��,�R	'��{�j$�@쬬`��;�僎�⑒6פ���I��>�r#7�ʩ��,w�qA6��|1bA�n��yQZ6�p�6�Y=u
ӻk�F�vc�v�ڔ�B��yh�6&>v�"(�]�	d�0q�(-�����\��D���E��&�P�k��bj�-�e�4�z�Yl�v?�>s/��{ �͛4�Α�jq77@�c��c��d���wO3�M}�g�?���K�0�Xle��{4��/�
�W���p�6�@hA#��ó̸���p��&�����N��n,�f�V\������w_X�DP�=�S�ϋ������ �J��'<��6�������I�yh����d�=v�|1|��&��WaP򱴺����� �mL�ߋp�t��h�[h��05�v+�L�����4t��cu
s=~��8��O�>>����)ūX6b���(�gw-u��G��#��V���#9�<�e�|몤ے�@�n�f$�QWJ!�KV����r��0�1û��E)Bq����ē�݃���=l����s4�����N,��}��̝@��l�FE@��$���38���x�=�m��'�W�g�V���o`�=w�ܯ^ĩ�<���_��M^Uk�SG��a��c��.��v��}u-�x���}2� �-l��t�z��˲r��)��k]K�.��d�ޞm�q��C:T.�n�Z���e�̷#w��ڛ��a����Ↄ�ß���36Nm��G�v�B6���c��;�ɜ�ٿ�vb��Y\U��h�` ϩ����O�L(����ϸJ�O�G��7�λ�b��2&o���Q�؅l��5�l#�3��D�X��Ǽ0�i�;�w]���c��ڍ4lAS:��-��Eg�L[���s*�@�e�ۆ1�ԙӡ3dt���5��x*�{l�Z�Ȥ���݇�C�E���K�}�iv���2�س^Zb�O!�^t�+���~�$ע��E��к5�����g���3��5K�:$𦚱�����#��"Y��s�s�-��E�h�_��v0閑��V��w["�B��ڻs?�?�~+
��3wՕ���?�/<�N6�i�u@�Ƿ����iYW.j������ɾ �G-O�y�5�kT�z��Ce+KG�_�C���7�i��w�h�d<Z�;�0��H,��b��qu���Xp�&�g*8�Cc�nu���嗪%��_cbcb�b%.����8��[��{(�H'8�	+����ƂҾ�s��w��{O�Ǟ�9��?��b]V3�lf2�X*�����X���1�0󦕖�5##͜Vq)�z񕠈'�̳�͋�V.��e��^�`\�3�a[o�Ǵ���#[9��꘽�N���8������N����������7��}ޮu��`+'N�YX��fQkY�>:�U�������r�C�ƺ~��U����9r#U�~�~���S6"|����e���y"�Y��F�y3�;���c��[Ea�R����sgpF��T��=���vmv�P2�#Vj�P��R�����@�6��	nq���V(ڤ3��p��c�װ�`\�WRu��zNL`�=���_���
f�$+�M����I��ᛷ��+p���g�$E��ո�3�5�+O�9��q��8�)%��UF|�
�a�3޿�c��T�i����͟����-{�a�2���
��o+П��o�zt�B�F��<c���}S�-���%�y�O推m��]�W�۫~�c�?�Q�"ܘ�*9wyz_���mT+A���HG3�
�e<�m-���Ae�K�5}��@0�mC)��c1����� ���*���Y�&6<�*���	���L7P�z'���
���Q\x�~�X>{�n�Sq��_~��~fR�W��_U!�z��m���������o�^'��(�@Ă�z�I�#C��Xb%��L��%T�l��Zw��Dn�`9Jr��Gk�Y�E�Pn;�]3�T�_���JPr���V�ю=���"�����3�~� &��L@�`g�rMR[�y����������ǰ]�`���oݬ�el����K��j�y���T]ך�.��P�5�Kp�=��5&�s��'
�|~��)̿�*�(`�w�q�^T���]���ʍ>8y!��b�{�RВ7�G��PA]m��m��������i����@�mq���֋���"�|i�N���8���WN�=P�9�ð���ү"�o}|��}+�*�b�gw�IO�R�gh��&��C�:�?�W��3?�j�C��I�ٸ���W��ɳ�Xf({��NX��,e�8w��]��qOQ�$��m���S?����c�?���b��{w����	2l˓��8�w7K�˞�n�*��C��ɺ+H%�\�����`�)�Y�:#k�?���15��̓?ƩÇ����0{�=pl�x� ���%��o�ο�[$�LMV19;��r�����;D�:�����_���Ͽ�_���?�L4���cxP,���%����p��	l*������F9�UQ~�Ֆ���>ސ4���5��jϊ\������.��{^�����(�d���q�B������ު�tf#ZA	��?v6�B�_�ۏR�*��}uc�B�3�S���m�Y�S����g��?�)������mD,�>��a�vFeMNf)d77����E>d[3qdO��ꮩQw:-�	 J�@ޟ�	�RF_@rui݅9���:�Coa�#��{�X��q�O"��!��`�׍�����m�8�ʹ(˾
}Q-K%Q8<�bPR��5�X�E��^<�B����:�v�R�,�2ׁ��pr#��߇3/������t(����X�|�m/�����&0�{ܷ��.A"S
hg�����E�篐��+m�7M����Uw�	�Ǳo}�.`���PdKԬ�_^�l�R>�vl8�/DI�^�u�u!�`�޸�S�+�)�3��r�� �������+�ݖ�lG�4O����^ƭ�"�[��.X3{��O�(���+8s����J"x=�"��˯¹g�{�5l`��v��}�Xk.��8�3������x��a��ҋ�N�P�oF��L����	Ο?���2�+�*�8˫���]�{��3>�����z�%D����@�dw���R|^���$N��:��]��Z��� �.�3L<�_�,��G�oC�Ա�C@�{�>�LJ��F4�y��^/C�9�lp	�҄��"+)�Z6|d�JUe3�x����_>����شy�C9@{����f��l�&@Y!Z��icǬS�Tj�f�!'-?)�c�\������$��x���\�Yݷ��Y��b��S_Z�V����Ⱥ&�ob�ƄvU��4㝽������Y�F.�]s�nז�Ex�xh����y�#J.]�&��'���h��~�>��yTd������ �W�	�s�}����R�1��n0R�:&y�	Uك��Et�e�[��ڃ�`���p=\�J���n܏�c�P�I�4��%���n��w�y�G�;_��Ls�Uc��>�Y|E������:�
���:�\"�i�;A��p�+U�ݺ)1�_P0ͳ��bl���wc�S�������I4�\k�[YH�Q�GsG���r0{�+�{�g8����t�3�y�!�S�u���ڳ����	6.�Œ ����Xxۯ:U���'h�WJ�zfU7B��^|�Y�w�������=w�[n��g����?��!$d��9WDhh�37Mz��xV�q�|X����F��v�mz�^!EA��YI_�_2�u*~s�&�-�f���U�=w�vdMQXVS�6Ւ/��Ǥ���ɶ�� �\[�hn9ɻlOz�4f��fg�X�.,ӭ߃�Ց�����Y�p�g�聒.��۞�,
D�+&��}�l)K�+UC�N'�>���d�U�f������� _0��5�<XM�f^�]Ξ�n���QL�@hvS��h�c >�<y�V��g,��3Q{�<_��a�����,���obBI�l\�1�w�4��V���^q�ɏ�SV#��37>V�$,dXEi{S46Na泷"z�`v2�K	�j�����s�,�/���+#�Š8q�,�F��9w�Y��qޒ��YjIֿz�K�4�:�
��Q�;E2v$��V�ݻ;�}���@�y��<pC�W������~I\�x�3l�i,�l�{��c4���gb�(���Q��ȸkD�&9�����C�GO����h�w;&��kN�`�歘�0����et����I,%�$Zy������ ���I�
ȠF5k�Q���W"�w�|'��C9qFw�F�&�]m��b�Į���R�����4�J�?֏������Am�:�"�g86R���h�%��FF�x�ǲXW=�0j��!cZ�,���kB�G�k�{vGQI�3�3�	��̱i���E�;�'O��J�ň(�n�G<6�pMir��k��d=��_2�4�PZys(�v؃Ʉ&��\��O�h=�ݴ=�kW�O�<�m��掔�"ȝ;�Rcބk7��_��6��}�]���]�x��GvO�8��*�߭�����1���&+����e���Ʈ�c[d�XC>k����\��Gcq����y?ڕ�D�x1���%��߷�'B��"��n=w��`	a�W�/��e�,�?� 6�؊-;w���_��˼��G�Y�d͚M��<^J��J�������X����c�?����ĭ8f�o�y�����t��*��I�鄦��&s��1�f�k�?�|xё-�Ȱ2���&֍+#�}fc�j�x��<���L������c���X��/1q��o��D�|3ѷ�Bo��rE 6�������,��w�п<�#b�7�.f�مz$`�m���o������_�k��'ؼ�z�z�x�GOb1�c��0���2#{�X�6WQ`�.d�sb3v3�=�2�8si��#X�6�e�����wL�N��YAS�U��� �:�)����<�R������{�2����*�xqA P4�1�Dn3�y��ss跺������:u�N�G�݂4����?Ф<s����Ҧ�6�]�d��'q�V3��}���=��N����3ՖH�Bn|G�$��u�0�6�ɕ�ױ�gi�����
0���5��$]k/�l�*��g�N��s��!=�q"�0zA>|QR�����>�3�±�~�zɇ��kvL����9�d��q���Kn��5��	P1ɴ<�(��~��<�Tnz#�)`���ᕝ"����
��������렜	 '@ؿ�P����'�0%�z��"�ԯ�E��83����(|��΋������^Ä��dٓ(�a6z��*�zs�Nca��i2^�I$k�T��n��w�h���� ?y��^+���\�a���dL�����{�~�GX��'���1Y��.��9�;����.g���d�L{{	qk-��F(h�e��i�.R���P�ej�]M\���}oJ��pU'����+H�/���a��!l}�axW]-B.Ķ�o��mw��y�&��qᕣ�Qp[:z���sM,Ûw�T��w_���/��m߉ݻ� ڱӟ�,��o@W,�7��/��\��c&�ņc��39���D(����S���dZ]5��C�y���*:�0	X",��C�g=o����i4�wUO�XL�Ru
�^���f�:w��-�k�3�M����d>Db,z�辥!d��ꩆՉ�o�<����kjY�"7�$���q�N�VQ,Ϥ�BYy�}���ض�e&/7ֹ�q6R�d<��댔C�_�R��Ry�E�^�z�e��@�n��nb��������3�L���{*hXU�{&�ݳ.x�ƺ��^��]i�Gg���ʈ6lö�<��GO�u�,�bfr�"Q�z�(T���ǹ��P��ĘԂ�&3׵����� ~T����T+
��0��
��5߯��K�����!Oi�5R���L�G^����S��0<��
n�qG�P�u>*�kH���.f����v��ã�2����n�9�= |�fԶlB��i��>�K�00�Rl�T�����X�3^�K͞���X�?����`?���}�!|�?���xc�?�����\�� ͽ K�/���m*՚^�g��k��c���ؿ3i��+��د/#H�9t.y��0Ϸq�h�`S{��o��*&�[}��tEb{�l�N�]�|T�d,�ŭ�ޤ�͹����u5�~�y|�/��Z��[o�AsI��� ���?��X��`啗0/VW����&���"fǶԶ�A7E�%X�"s��MB�s�R)6ѕ,H|D$]�N�K��}*'��6Rk��9������� L�B5��K;�f �^��zH��R�n�~?V�}�r�� e9(���kT���v�v��"�4���EdC%��kJ�B�L �Z�W�X�b3�y>L�`���q�Fq/�D����
(���[>�b�k�{��I��G��.�$-Ƈd�#)RO�b���������[8���X�"8���Q`�
�2�Q	�e�c-ny�������سw/z��yP���q9d�"?���	�#)��S���΍���XK�]��?�9^nڣI�\��<S_�,�;nA>]E絷p�ǿąwO��e;�E�Z�ۘ�ڌ(�����]\@%���7N��d;5�KO"�0Zw����s���?g��D[�R�L�4������I���Ҕ�h-5a@c��G<�c��}ƕ�0��_k�Xu�$�ؕa�X�=�VO�{s瑞9�� {Sn�mR6���9���(�܃���q��؋O?�A��C�{
/9��T��g���݂X��@ �+��%]4�ډ;���x���qv���Q���������#��ׂ���:E��h��!����X ��i��*��H�1@O e���l�(K��t���	CO�Q��nd�?^�Q��&3m=���M��|����k/b���R/F��A'B�;Юn,Ъ�"B�I����u(�jf-*'&��
s�KgXU0J���aV�p����剺�3v��2cܱ�i͒d�F>��`-��G�'sa�`�}.{M��M�ݍ7_~s��a[���ܢv���	ß���5Ͼua�--��iF�X�������q$�J`��!����<>/�.�3��>ڝ�DF*b����-��4�ǲ���$�9�:�3�bw��E~�G|�c�1��n:��s?F�����_���������Џ�~_AI�R���p���������/���^G���u^
�Fk��}�|��b}|���sT�G�c9pA��$��?H�
�f��Ccc��5�e]�[���p���`�`��:���r�t��r�ɬ�k��������_��;o���+��z6�`ņ���7>�0��j��D�w�|a	{fw��_���m��O�����A*�7]�q��n�fw5�]{N͢���T|b�W�sc�3��_(tKCZ0��c���B�E���'��bǘ�Lf��>�<Q Ă[��^��7���-SN]�ǩ�1!P.�vI/�=Q4VUa��۔��V�����N������D*e^e�z[	��*�IRC�z�Nu3˃�o�����h��Ya�p�mg8���?C�q��<��0�_�^CfB1�R���~�`s�._*���Q�&%j��y�5��#�z?f��>��|X����s&���W�~��U��qmށk#K��h��;�.d�u�$F��x��9:j=�<'�Nq܇�Nm9_ʐG��1au�V$��fk_�&�R��0	�#o̚��) {~�Ϲ��� v��g�z�U�����:*~�J��^�p�oD��g1?�B��`ʯce�� O���y������l��c�_o���:�̡Vm�]�� M��4}8t�}��{դ�U>JY��fR!$�K �2Bv���#Z���O��7yf����u�PE@�$����(�Km���3�{�e��a�g������X.Ƙ{�=~��|�nی���������5$�1�[�$R�21H4��+	�_��s�b��Ey�- �'��%�7B�L�v��N]������y\(�$;�2��6�:��Q	�^������=����7lTv>M��p����Eb�ڄㅱ�fB�&K����(��n���,�������D%���b9���['ى.ײ!���<T�@ױJ�n�"��Xu{�f�k�S>2<1��˰Є�b���%9�s��wVe�y��	/9E�k-�1���R�QL2���'0q� ��^��7���e��Y�n�-�^�Pf���Z�]3�-'�fto��F|��!k
B���V�첮�B+�hgQ#K���������L�.t�JXn	�= ��̵"�R.1]�g�荦3��Ow�v�+Z��*{�o�9n�͔ȜV�«6b�ȃ��e��VK�|�g���o�[�!�l�X^��t0�X�t���O37N�A�.�y��O<�/����>>�X�1��ˏibT>`�������4ǃS�ל"�Q���ʹ���k�P6�����q���^���$/d��N�Eʁc_����^� :ID�]�X�,��	p���ߣ%�]��VL<� ���`�숈�hb������ܽy���tD�f65BX˜�,��j�I��4E��e�M�s����KM�sLPv����D ��ȣ<n��i.֞ ��O]�k�\�d/ڲ��50=9��]�c���jC8@������{�ҚW�?�#Ҷ���*t��!��&q����w��7�ƀ4��i|�>�ve�z����ƚ�NF9��5_@�s��W�8PMRaf3�!Q6�]>nΩ2`+���gýS�W�E۠�j;5��~�����%�k,EE����!��0*�j��؅#g��Ⱦt�,��l>��mV��9��럂�쯉�	��n��j��^��AM*^�P����l�\	ɾ��B%�Q��+�"f��#?��S�Il�']IZ��8��*�Y�ź}䙽�������ܘ�1����ف�W��]��x�U�Z���b�p�8�r/U����yL���&��=/���J�E�?���ϰ���0�u+�c�u@�C�(H�nO��<�C}���^��t�Z��+\����Ja��7����!p��t.���1�
�6�	?#K����&��}o_a�V�5*�s�=�=ss�����D���ؽ��w���}E����z�T-m��&��B��5�1��/\Pf4v�+��-�]ގC��`���L2�0M�W�p\n��r���X2Ȟ񖞕�v$qɜ���S��۴�>�0���X�E�z[�Ef���7?d�Ks�g�`ڕ�6�o�أ�$�.Э��rjߵ����?����p��Pg=����]�j�H[.V[m}.�A�\�X��Z֖�}�Ϭ���6cV������N�S�!{��/�q*�Z�`J����k�$���ЋD����NԜ݌��P@K�<���
R>�ĸb�<r� �b�Y!];δ$��\��~'�7�b�$@\�{I,ِ��;G�<�����W�2��Zz���Z&�g�Z-D)������n4�J��d�Ej��p9}D��M�.���}�і�iS����(u�6i�E��i؅��Bb(�MW;͙ͲQ���\�aj�%�|я�>��紆
�v ̭��q͚d���E3�-��mB]�~�K���_��{��<��I��(`~+Aؘ�+��.0Y�6Oz_���e��C^��{\���|�1|��׭�2��#�o}�qMs�X���f�ݫ����~�ZD�Ɣ��J5����!/4��Gu��o����n�����^�lM���m6���a�u��V�]z��Z�x0�h�)dw�e _�=�i�D�v;���*N,�G������A���S/#a��k�}*?t��<:q4sI�vWp�'?2}������w�l�8O+E$Եp��F6>a�����^�Z�K4{%W�9�o�{��뱹��P'��T��^����E�gz��UdJhmZ��i?Q���ұ��c�B��7_3'�ʍ�b"�Wڳ�����?���K�+hN4���l~��եE��Y���&���Sf.QT��ֳ����3-z�,�����-�5V�;�U_���N�*>���j�+�]^� �6q�;@�2�����.�p�0�d�☻�1 C⓮̥1�|�����w�Jt/�Y�n(os�u�G��l����N���6τ/
�|  �8����BF��֪R�2��u��I>w>����hEsC�bȊzT*��d�q����t��59/�����Gڐ�
9�;e,�l�����n����z���0����
0/H��4*�Ό|N���(Y54Qz�86�7��#��r�CVM07XA�D�����	yFshV�Ι$�����s痲�'|�KY'����G���h%��"X��8��l�=�a�$��&�iL,3聾�� ��$�1n� ��虒̠���W���\?�m&�:��'�r�{p����r�G]ݼ[g����P,��N�@��N�}��n��C�ÿ�jN�JԴ9u�I�K��Ēvg�|���?�9wNc�i���A����G'�z6�5KH&��CW���s�b#�4�c�Tl�:�ag����e\�q����z�ܩ�ᘙ0�4��L�֔�y����1F�Z�6���`r��t���j]qN�W_�;�ſ��ݻ���c��{XK=`��K&��_w�*�FweW��t�F�"̈eZuCuy��GeG�Sf�-,��g���e���`X�l6�Ec��Zj�DÁ(�m����J�Qא��m�#�0��a�!�d~I��v�}�8�$��(�xJ�ބg�cR��!̵dV����$:i�{�� �'��ƅ@xec�T�bU2����;S�a;܏���3���_Z� �O� ��Ԫ�z=���lr*�����c�CM�72��W����8�3�%���6F>�ўٸ�kc�������+��W?��o/`�g�E��)��䮍�v6DAi#_ma����}4�>ʓM����,��ɕ��M�{s��L�d	�6���J��u+�C�u@��[_{Bۅ2Y%��Gi~�S�+��@/��SC�c�&�6umv�cK��R�W-,���=.,ƭL�ߒm�x�H�9Wt��R�^$�[wY��Z�5��⛖�T����Xc�aܘ]����U6�����F���7Q~�^L�s�M��%3K���$��w��o��Gv�=�x$�����C�_]��:�U<麥jU���m������-Z82�����r����\@=en!E�/TB���C���DLO9�Ţ
�@�l
X� ]�dSP6d�|+���y����$�U0���[�U�9�j7v�|������?�c����%�)\#$_:���%������"����ާ+9&��XC�c��TA���yb��q�!���3[,T���	@:��hK֤S��߽;o�3wݏljZ��Pk۝a��n؏ѣ|�Y:Y��g^��ql�e���;oǙ�~#��!4���o6J�m��[p����D����'V.s��(�������C�%���R��*�@j���/�s+�bƲ�^�+2��ʄf��9�E�>ϟܔ�qwL9��gs�Q�;�}�] � �T�q�'�6R�s�}�܉�3�g�ç0wb�i���X������1}��@-��s����yLt�PE �8���qLU���N?:�/Dl�k��<��a}|���r|�+�k�5�O#��0������"�:٠�P5|�uڹ��L��U��'³4��rn5�<�?��Y��a\��;0��#KM��u���3���I���38y�pǶ��##��D[�����|G.��Ɉ��_<`�o��[o�̳�a�ΛE�ߎ��qe��<^y��8��g�8�-�rY������9&��9薝���)UV���nf�Ԁ�L��bX�lS�<ka �ٌ�ߔ�uN.�����q��@�F#���K�0�lv�p�ĩm�B��P�س�Ťxd�&�)��f+hv|"s�f��y����N��0���f?����C�0����I�J�vy.��n��p��B����Y�yW�s��)lq���AE�mY�j�4����8F��g��Ԙ�/ ݕ�+�RFuzuЛ���-�#ܶ�4��EL��,(���CU��c�c�A�d�[*T�Ѽ�t��c��tӵ�p�]8}�8��U�O�,2K5� ӵ5
��������2��Z��;�s��Yi�b�R���|�B'O<-j�/��g����O�"�m��gٴ�+`N�%�F��nr/�RI�.=4$�n�1`�s�������F�����yT��J�c��ITj={�m�����>���V�6�sfy��%;�"�ވ�l�� �w:<���
�^W�_�^�� <���p�V�[�*Oɾʘ���/?����>>x��������&.ʲ��>���{7�b�--�-�j�hl��J��"��ò�\m��;�����-�v(�� ��9{9
橋��8LL�`�ђ"Hz&��������k�^a�h��/����\L5=�r�(G�i�]Y�$*��!N��*N��&��G�7bi�h�]���74�
zb�:"@+��]c�GT>D�b�k���[ǲt$^�4�.A�r��1���B7,�?��N�&!%y�EQGf�n�m�=�Ҧ�"�T)�"������)��rz �u�5���)(�[��A��X8��h��F�*f~Pհ�2[�:&��Q*��So�u-�D������u*�P A!w��w����+-L���]X�#
����p�W�dmEys��L��Cn|Y��=�pGng�nމiT�l�ԆM�Ln�Į�pw�ۨ oVds�ςP�^�h��l8�>�ٸ��g�I�w����*����Ŗ{����~�X�tzsؽ�DO,#�����&2ӝ�lV�l������ɞ�7�%��	�rm	�z;VA�m~.U&��ޅr'd��hYe(�@��Z�����X�A]����� �G��UynAI�a�Z�·jU��3o�p�U�.O�>
C�!��_�輕�ׇτ���3W!�<�h�x�O��|���yo�_�w�����ϣ��Q�W�]^����]q�}#��Wc�=��r Ϡ\�_<�(��?� ����:���_}�(�b����Q�^���?�Ԝ�VY�l���n�4�����M�c���l<�����1�Q�j�s8���s�H�2i'VZP�4��Z����r}[k>Wlq��((@h�P�S���D�U�,iv�7t�2^�%�U	L�-&����ˬ���g3^�~�v]��r�Y�VG |p�^v�hܻ�� j�d$��)L�ј��j4���cH6<uu�N`�j��ێ��0�]��iK�VX&�0��|�"�wm���`�m���o��E����d�d�sa2����$���}3�.ԡ��[PS�,,'E����NhU(����OĤ梱t�,���պeC�f�B���Ӽ������K�:���6�,�q��6f��"���L�i��,�;o<3�O`�9��`FKp�^�䖭���L͘�3�M (g� ��oc�=U������p>��ڕG���Њ�W��t��-���!�7����a��1L�Y�Y���&,�@7Dw���̝"�D�
*�I/K�ߕvKKK��MֳZ� ��]���"��L���=�Hq��欽��p��@���΍�*�����Μq��T����")�^0�2�f*el� [4L3R'FPq�si>��_T X�Y=ێ��Z�<��L���y�	8{ ��,c�S��){ϝAv���*�ZI�TO�������S���}e��c�{�T��^��/�v�ΔKE.}W̗>K�偡�X<��Cj�.�.؏9G]��C���9�kGy�A�jBK�"3�܌�j&�j�]�wߔ��bx��Lpf��1��ZBL�),Cf��=J��^}���g[3f�+����kC͒��V�>->��0�&c&z��̽&�a(���ؘ�2��HS\��T<X���}�&*�KY�N4�[|�{�ܐ�8�ٱ�a^7Lr��%�гX�Io`z���v���c(K����Vu*��yэ�!��V=T�lT��`���L[�J.J�e�r� �� �qZ'qj�_�cR]�V��&�PmT�+=M�R-�%S����&5����k̄Ƣ��j�#e�/�����r>b5��^�'�MV�=V����$r��{f4�=��`�F�p���� ���H�Tm��:Fpd6[�?�c
M���z�����7��0�
C\zv�\�\�uʚ��y�-8���E��* ��m�0�J&9*��7�{��DY�m[٠Z�DO��պ��y���J3�]�V�K�KG�L
��W��r�[w�zuD���U���]�n�� �(�S�qu�̙�a=Z�������L��ɘ�2a�^b��u���4�!w=L��&�Hl�K�<�*��.T���j�R?�
d/�\�z�f�S�-���j�юI�����#�{��>��(���9��w���!�����<�Ҟ(��r0Te~�%��[�Y�%Ϗ^��+�[��<��/>���{�	r�7���7���]�Xe"��(ͯN���Ju��n��)'SQ=�,��"�Q9�i(5�V�f"�c�Bi5Q��; +Wl \�zW�ھ^�I�O�;��5q,7�"iaj�++����tj.�6�[&�{ʉ4��;5~���~	�ȴ6վ�Y:�WG�˜�T�.�&;�*3
��pB�Ak�s��c��R�#�9,�):`壤�+�\4r2�5%@N�u觘ܺ3{��%���<5m-���b��K3����S�
��[�̜a�l#��kIE 3>��v*�wy�uh���J."�dh�]���W�$+íه|��1�t�7�$����i���9�Φ`�s̜���p�G�C/��~�ð*�c^��M\�t����yjf�;rA�N'���vΙ����l�I�+P������1���M���ceX�n�t��}�En�kc�k�"���X���.�d�3�u��NP�X(f����!�eD?N���D�v:�ːj�Cn^C^�e��6S����8���_d�1�Mٙ�^���G�#�����Q�1毡	:ɬL�����3�A�e�^������g~�^���͘{�u,��:f��n���7qz2�ٓ߬��Y���k��g�O�����d��n��X�J�ȮO�IGIV�vP�[&dF��9^$�����E7���G�&H�F�g����>�`�e���%L��Kb[�a'�jWc'Oз�v�y�Ҹ�,`������`vj�����Z��c/�\K�B�����	n3�5�VϔzLvK���K&��b�IӮ$�����K;3���3HaX�(�{����Q�O:�k[}���v�Zc�o�RGs�f8ղX;&�̚n����[j�X�;��*��\ו�1�{�\���AAȑ��ѝ���!�>�p��0<�fe�;wIajj����<�{�u�J3��@&qQtl-u�pY,�m=���C3G2�)zR�s��=�YU��fȂ঺��-k}$�Q�Ԅ��ϭ�c�"I�`�5�~O��<&��n�J����U��B/�=��g�+��3J�� �_udO1�OB�eM�d����g��"7��iHe_�$���З��E��-+ �c[�,.\�5�}\��kL��Z��~��9v�a����\0<�IQ͎~��54�w<ɳH��ͺ��>��o����(��S�O�����P�)jB���2��1���M��
Y k�qQ��@4ՠ���+��Y��0s^LR��`*Zo*�Ϳ���������:��������lG�KװWJ�[D����T�y��b��T#�@^X>�*ͬ�:�ML���3��5�Y<��:���cu7���M,d�&SX�fL�됬g��@?��-^�%I7�f�G�k�Q�WV#�;w7�t���j�쩧�6W�����E�XI4�PNsI�����A�Œh�"p��ճ�c���]�X��M�)bv0Vr��f������#��+JУ���ռA�C76���G�*H0�ͤz�)<�c�2iE��Kb��6�����f�69/�ԋ�����F��4�N��p��q�۹�zr_�b�xd��ϡc(O� ^�
%˱�G1��r���Q��L��o82�<�R ψ�y��u�j΄�ld(��.ϒ�i*8��I|D�6��'&'���æ��k-�"�l�����%�ET� �ᤋ����w�<�{�5K_�WE�D�v֢{��r�n�-�Z�ِ2B�P��H�,Z��o	ȯ�^Mh$��x�2����Ԥzsί,�L�o��zwh�3���py_5��sLF����	贾C�6Z̎����W�3T��a�0�e��"7�DÆ��[i_;�HE_	DN�˞�-��(U)Uԝs��f.NL���#G��V��T�aT�C�����y��|�Z��՚A�~-�g�o}/�M�G���dGq����dI� +�lɏޗ�u�dQK��c�K�@7���^�zo�E���6-4�a^�_*�6=��j��*����Yv,��$!�s��+��*���cCl���VpF�bI7q�Q�M!J�����Dy���k����gLʽ�s��^a�*.�n�aԽ� ѣfHr�(V¡G㒑_���7L,8W s�x��Yȵ�W�-�`�[�K��o�Q��e�����Ӎ��$^ճ� 8#p�򹓏���o�0[�\�OxD2�lG�o�;)�BA r�݂���Mۤ���;ZԳQR�?V=�1��>ٰ���;�B̭��J��͑hh�������u�\�a/@U���k�#� ׍^vtJP��&�v;�\���f��Rt��tH��1tnX����ߒ	%W�[X�<a\}�X�̡-��&}���2��5��k"�\�;	:��5�GL+^5�F��cϵ��/����ض�0aC�j�[@EG����m�AA�!S9�9�Ҡ���%��<&�Z������sIz$��{h���홬m{�h��>�c�Y�
�Os؍���m�3�VK����z�BM�<){�Ka��P��%�'�mp�����X�+����5��\Eu�<�~��~tGT/�x�D�lc�9�2w�w�Ԙ]9 r���HW�֣���4-��uj�m9D�rЖ��oѕX4;��Ln�Ecj
ac
A}RKsVEkA�kW~n���r�؈��{��V�b�Rǌ ��r�����շU�=w�<�_X�7`qnI���fQ�r�r�����֪f�O�JX�F.�VYY!����f+.3tCKWY���q_�wN���$�9��}ma�'���d�4ft�Q�E��M|�����r`z�kݛWl�o�w�0��p��Ė��~C\�ǔSӪ����<�\����'@A#��J�)	�ibW�&s�f+��g:4��Y�}���Lg�gQLf��E� >��=�ˁ~��?`qivH�d��i��nAƔg�p��)5��K�	a� O��,�B�X��ns/�0D"�zBX�g���|�0w ���]�U��8��nn�uʥ���!d���;S���6}Q�:�ZG�������rI^	&��� ]���G�*�QN.[*�0�%'z�]�ݤ��Y����&�ZU��פ��Xż�V���3�N�Iy4S�K����e\8ss�0�uTъDj�|4��V���4�)�����!JY]�)�V��4�Tm�����Q��e����c�Tㆿ��q��F�<��ٛ��tH��&>��o|���}��ұ���˟7�D����F�����NB�o)6Mvp�`��lb�\Ѱ�F��,F,�pW4�X�"kN`E�v�m���>��Әܶ7^s5�F�X߾؞�'O��w0��%��%6�nG�\�����&�s�D���E5,+�Ĳo�kh�ue!�ٱ[���rh[r��jK~����xf�S�,��ߒ{Zm�!7�`FkN�_��\�����k��Z����[P]��|�L�X��?S�	�g7]��n%�����3��Z��5��0���}펙g����mk�a��
&�LAB2��jL��a��ꂋ�r6�N�PZ��$���C�Ze�6����TǴ	l6��H�Bfa*7ɁE�E�-0MNQ�8������о�)�Hw��ڿ7sP����7�tC'��z,̡-_%�1+�_OK�����&��K&6m�J��ou=[eh���,sJ&�J����q�cd���)�踾��8<��f'72�s���GO��SO��(�ƥ�bI�^=vT�łe�ۆM�1�y�X�e��vDQ_Pz�	SSӲ��p�m]��4eĊ����ϩG,t��A����
.�j$�o�4��7!F��I�wc�M3��`%ϲ �ܙ�8y�8Ο=��s'pvy��$�3.6Vj��=��u�Ϻ xI֣'���چ�J�KD�V �X:�à�G��@-��=`�Au)N����r�M*�i��y)������%c�/3X��<�/`��~�'�<<���}an��RR�>��F<ܨ��̓���ֽJ��z�dS���YO�%��l�-7߂�7߄��]��S'N�ͣ���^Ù籴Ғ��ƊX�4�C݃E��1-,}��64��õD��ɧB�IA����R59@Ur��\lݰ�H�}9č�인��2�9�.����oFj���m'�8O�}�E��d-&Dx�,�.��(-��E�~e�Z��eK�.^͠��ûȳ[ �����������&!��q���-�>�x���%'W:����0u�z������L���F�&;���x���mj�?��,+�hE��ża�O�����8�<D�,h|�v�#����B?Y���s�+c�2ȭnw�g;I�j���h��X��ѣ螿 
,s M�c-u*+$?ah�!+�pS��<�\3��`lG�,mZ�e�3�z��xR�آh��3�J��ٮ��,��GZ���N6_���Ŋ��{2����gђ�nܺ�o�����{/���L�{�rUW�FND H $A���$*Xi$˒%y$ٖw<�7���'vw��9�Y�+�#Y�,˲I��@�"�st�������������=g����]����������.�c�-6�%�=�d��(F�G�q���cV�qsꒊ�-�"�jkm��CK������xa@4QPW�o S�L��+܏�1��X��kq���� x�&&��ùKgp���%��gY�a���(��$�ٷ<��q4sS��`�3���Z�ª%=�Tџp�+~kw�
>��՘o5y�M��XO/�}���]����_~�#���=�^`%;ބ��|��M���N���$N~b]�M�&��5ED�4Nr���� \Yx5qp�‹i��ˀl�{|;��GM��)����x��I�^X�h������2]2�\~�ZM���t�coR�P2Sg���J�����9�DK��a�&(�*_���3�9\#��@�fI��f�ib�=� 6�Y�u�S��(�Ė�bT����c�����u�ZiqY9����ug�{˾֮v��z�N� ���~�:D�������K������m��U�f��D��>�D�_K,>[������(��0����:Cg�y��SK��i���`���* �W~A�:a2ۊ�l��0���9Ya���!���2��m���qY���fXS�EoEt�������w��{E݂�Wo���Y2�,Q>s	�ݰ����J>\5$8u��B���o�a R%x�� �[�t"i�2ˈ�X�{5]n��N�=U?�\D�m�,�ZP���8��|vM�OU�2�4UyN�
����\/R�����R��[���V0a��$�/u,��8�
�g�$�]G��T\��t.��;طLZȰ�I��-��M$U�`�w?`{\��ج��U��|C.�5�)�ct�����=w��O��zW�^��W^�ًWqY���X&�c��]+�nՕsS�[*T��#�6�[�p����s��t [�L���1�~-h�^�j���7>�)|��w_+�w�;^q�t�P��1K��)�G��{^*�}���+�܍i:�/��ي���L����e��0�l*o`l�.<~�A��\G��'��7q��e,W��D�(���d�XBG)2%�:�D��ic�M�X�*�P�\ӹ���7o�#��Vw`��J2��'�z+����s٬f�87?�S�&�s6� R  ��IDAT�fl[���kP��Cea� ��C*����B�)F*�##V!'�4O� %'�; F4�6��'"c��ft(��z8D��
�"�P����.G���|���t��g�X�xg.�߀LL~��ҳJB�xg�$L��8�U��1���+�fQLm6�U�zD�R�_�o���
���p8����+�?�������јc�}���vh��o,xн뗝�;^��o�g��_�Z�+Z���6��6�N���u%x�n��ҩ��b�u�f�ު��5�c�B)��[��M�]��mT������F�ӥA����_,��R�F��k�]}�$���֑#�%���dո�e2��I/��)r�[� GGT��!v���<�-A�$l�3�?W�b�ZBI�-1�4���)��x��5��8\/,�EY#���� O�c�� �ADڞN�-O!�
���e	�
r�/ߜě'�#/H}ˮ��{`�:���?���2N����uG�g1* g���n?��R��U���J'�>�� )[[����"�rKv4j�ϻV�o9Ӯ���tۻ����u�^��5�"�\v�c�K�;��&�;˕��C|��1�,�mR�A �r�@SP_~t ��>Td�,�樰ּm޻��Ll�eA�?��x���8{ZY�|^6c�څ�l�l:�v�-ȿ��j).�D��������g g��_���'t$d�J���1V��5	h��Y"`��J�U��7�$��^S��W0s�(N]���#�c�����-$�D�i���f�p[@Z�	�9�Z���͗�����J���%NXI}�N�wa����alW	L9��C֑`�.�7��~7�-[����+Q+�Xav;X��������9��k�D<ʚ^}��ʱ�_��ö�n�>�U4Tŋ����a���@%@|���A6��m��SѺ�cu�覑:���_z���o8?
��6�>��+����|�40=M�F3�~�Z�"�"�P?�7�a���v8�Պ���K'����Z]	��� ü7b��Nm0 �;��,���5	��$�1�-��-��*�k��7� ?���[�cz���(����YT�!��!3>�m�3ˋ�.-������/N��p��U�	�Giฎ�uU��N>��5�0ȌhSr1�l�p�L���!��k�&�"E$��!�?�Ry??r'ΟGV����މ}{�b��Ob���b��I�{�%\^�Š�cS���h^>���2ҭ ynɊ� @�"�j��U,@�S�^�`����X�C��i������o}����Ż/�zס�z�����O��<����b�{�rn4�t8�o��h�P���vb��!�*z0լa����];��ǐ������w��#GO`r�:h�=9�$Rg��}�$�iP6gV��B6��P� �=Y��=,�(�#�
%�Q�T4�GbKJc2�E���t-�u��k��E����f��3��ZU��� qS���$^�üDÅ�[��0��D��0�i+lA���(���}�PM�4���q��Ӭ+Q��O�����]��`�*r�Q�7*��W��.�M��gj���&�&�&#�6u����H��UR4F'��+�r*V�T-%�YF����i'S=�PQN��I��������/%����n��H��w7�j��|�,?��w�]�N�j��Y�r�+��:������F�(n���*�G�����n����S�|����+
s������}�c�z�Q��/+t�ijȂ��a��K�+~��1�yȞo�E�I�%�&*r�	���^�@z��BM��{00�F��ƹk�P)������f�54��k^����]1�t\�Qxl7"A)���S�̓)Bڭ�NlK�Rz(�=nNps�P�+���j7Q�,mM J��� w�A�ҵD4o�����T�y'��͸X*��W����3زe<� ;���ۇ�o���G����4�l��1�r-�4ˆ,�d��,��xKlG��Y�������-����&8�7�û��׻=|��'>lF��c�{m;�`�r���}�=��:�);G�鰸�LweSp�H�Ȇ�đW�b�}�a��p��4��ַ����]��3-F=i]�����(G���x�fxkFǑ�%�e�Y������<�r~m�\_A� L��Pǹe�����ڂ�ҿi�9qʫ�� ��V�^���("�H��W+�^\���;���/0���¤��5�<�����`���bc~��Zڻj�����p5�NX�D�|B3
����,V��M�{���]��_�g~aH�*Tl���1E�L���O ߐ �1�m+�=;�$TM�ba�?L���V�����!���,��ֵcL[�:3��_JƲC���D�d����w^�k�
�XǷ4ˠ������C
��FMtZM�=��uk����l/@4�C�nt���Z%�����_�������xƖ�-���}q8�\)f�?�R�8X��̛o�r���![U6��`�ú��@XBn���!�C�]�J���� ���wW�y�-FHU~ױV���*�]go�(UkQO���<�e�����N`N���r���}�=$x�qkS�� ��3: hA�)����6����:�:[VY�� �t�r�|6g���6�٬��j��<ʈ����u�#�s��7���O���e9G*M2��3ܩg��Z�b-���%j��x�.%�i,�J8r�,�ݸ��_�9�8x=�l{�a�}�\8�n�g�޺����_�`bY9�bE@�R]�bI$e�UY������Ŝ�B�)gR��� 寿�Y|���Ļ�wz��#R�(�0�y����X���;!K=#�+�f�c���T��$�ݴ��u�{���������Ǣ,��z	��g03��ӽr霢�Z���,Z_g�;�ȏ`�����'đ�d3̋���u�gft"��6���Pi�ZM3�������儒�)��K9���6�5�\�p&�)��[U�0'?�d2H�Қ��b��\T��Nl�Jq��I�7�%	r+���B���3y�b��A�e	BZr1�r�r�E1�bD�89p�@"g�v�"d�q6��OK^�WyF}���#2[T�6�]չ��ig��f4�d�{iS�~#��H>�O���W۞���0�o� +��a�Ug�s K{�y	[��v�Ӛ���s�y���5j@Aj��
/$�G��3��α���c��Fi��H~v̘�qN��b�AP�%�%�	�4[�v��Z�31����lG��PC+��QM6Ծ1�J"�?l_�:Z�����^	hI�r�q&�\\��S�ZȦ(�[�73��������C@�}2hVh���=\$��s�b�~:��h�\e}y/2����N�h����Ho��V�fp��Q4n̠u�F�1��Qu�����FBՒ��G^��0/�z�R� d_-&m�j�x���1�i=��;���N�D�'2(˳�ɀ�f%x/���N%Z=uԜ 焄Ru�,��6�Be�Crd��"a�����{�(\������GB+�CeI��#O&��O�%(��%qy�G�	�A�P����=�6޺t/?�}���cO�����x��$6�2ؼwZ÷0ssJ�p3� �ciՃg�cL>T���k?����-td}P�����ݗy�������~R�OTG�l%���Z���!�MpL%{D)�!�n�j�,�ehl��Q����Z3��8��7����Ǐ��˯���"�b�&�m�Q��Rłlhq�I1��w�ݳ{��g�E�X�ٳ�p��ܼ}Ku��v*.N�Ӛ�����7�JT�8���B�Uˌ4Նzn\
�D]K�t�`_հnɦ-�
�f�'9��	k�*!�$�F���b���}�v`��X�}S�SȤ�J,+5�(�c�������jj�t.4ۉ�`��a�fF}9���o��1���ê��ʫ�4W�b�Χ��#�n{�
�0�R�`��AEmqꂠ< +#K>g�vK���s�ՙ;a�x��H@���+B�	ZT#{q[����h�=�g�p�tچ_��/�%���|+�yazFo���8+e�Za�p28����A�m�m���bfX��Co4O	
A��dm{�	e}�!�-a&�PI��w�+S0*l�3ZIt9�X=�4Pq�i�5���a)1yN����+�?�<��:���e�7�Ѩ�����wF��D^v(�k+I�*�0��}�w/Z�#X�J $�6�a+��X7��|���:}N�zi������4�e: �ۥ*�pI��"y$�K�8ݹZ}k7���A	�g��K��P�!�?O�vA��"��*�ݐ{Ќ���H��p1$��v\D�����t���k�n?�
[(?lb���uѐ ��G	qf��O���������xZ�-�����9��XA�lM�M,�7�>3�KS?��Sg������q��Q\9�:N�yl�=i/^AsQ@�g�C��&�OO��.t:�&;?q<�E[�W�TF\��7~����_�5��׻P'";6G�z~�񽧪��ƾD�
8�H���a�%�H� �~-�ܱ�׮Ezh%�8����'���iA���c����0���K��%�45������q�=bd;���Ù�Ӹx�"L*PA,��Z��tMe��=שPa�ԋ�u�b'f0�����o�:�Q[�;��=��׋ڞ�1C�q̼�?��	9.�)'������wV���kp��8f������b�im8LʽnT0�Lh����Ũ$\�oj�AT7���;$aW�V+�X�S�0?�M�3Q��
��V�L��v�♳gQoV�/�?��#�M������/�i�Oz��c�Z9{[ۥ�0��^l=�T׌`���o�U:Z�s�f�����F%K��B�c��Wn��{.I~4�ay"2�R͚.���U*ㄭ�G�k�^Pÿ;�EQ�I��<r��S�������hU�Tk�wk��Z�;+1�$4 �U��G�lsY_��q��gм|=�
N�L���� v�oJb�^���d�zi0������[P� �0}���Ѕ��Nwn��g>�k�n��ѓ���3h�ej�[��3�P-��cS�o��{��{��k�~��!\�:�_{��!�n���8��R	J�&%�4\�IE�t6����FHh��U`�z?���5��x��o�e�
�UD:��}���4�b��E�B{����c�����g�`W����kՒ��j�*�Rb'7
�ٷ��?�����.��מ~
��#3~�>�O�<wkd�M������XU�:z�k����l����:�ǚ�<���w�_��g��}w��v���O ������n��wU��'�f�T�j��ˆj�B9�"%�<�i�~��$�O�h�ٷ��\���Ėm�֛��V��ԉ޼r�D|��p��$���8�W��*2P� �)��!.6G�!�4��]r���nZ�"╦�C�;�u�z�c�����w맫6u<WT�L�f�8=�HN�1K�W,���albccch�
x���$�x�㏣w|B7�G-hAi�RQш9瘢Ϡ��!(���M��N�ӷ�q]a��̉G�>:���Фw��X)�F�$�LMvϙ�)�nb�[B�D��u�
(\���mwap�N�$p�'�8
Ӱ�͎>$D�I�넁�9?+�X��mN�n�%ɉt�`�$%�;Uy�$�P:$�hhD �qt,��u��Db&mC�J���[m��{��F�\��l�M�ry<J��!��m>73���	�1����*�f]�N�Z��ߖdGު鰠`i	�s�Q�q���gv��2�N�I��}m�L�{�K�Y��Q�}���\�텻�\>q����]��ݐ�@�XZ���/���?��O>����#��҉S�s����w�#o7Tt�*�R� �Fbh*��%�8�^�'x��˸1;��[w!#v���+��TF���׼�ʠ��Sɖ�[�h[�٪���%;+�|7�̤��a��.�n�w�yn8�]���B���r�(���vx^���C��y�:wU���5P�^�-^�X\�΄>�O~��x������/����q��9|������~���������f�6��<n�>����a��V��T��R���Ob��l�:�jn��\&�;�u�:���7M������#��C�	>f��kD�~�ـ'�|^�7<wt��[�a���q�~x�>���ï��D��%
ߵw^y��_�BqiY��w���x���r��\����i��5�E��L��Z��1�^�8�N#@�Lvfs�v'����^���k��7�em,�����T{���2�b���i�N�>�^�*Ku�a��_*,᭣G�s��{7&�����8,�p���oێ�[�5sA��Is�$i�1l�	���u�#3���/��@u�����Z��a9 �������ל�M@�<Vyvtl�7���-$�ٍ���Zû<5���Gk|��!4c$�Ȯ��]�5�#S׊*���D<�����r���'��J���TW���g�&�SJ��䚤pm�r>���$ىx��D� k���X�v��ZV�H�����#F4�5Ȫ���~~ϴ.vx<�dٽ�j�P�;������^{{�g��U#�g�W?k�yw�F+ߏ�!��<7N��j
��ʚnШ �S�:y��@��Ozd�Pő�<3ߞ�.��_(��s/�xD��L��?��z��
�~�=��q�a���'?�qAԏ���q:wO|�3��u���e/4�b[��Òܿ�S�s�gU����"�����G��������ؙm�@���gQ�{2�m��_���B����aJ�P4���@�;�!r�x���RK,�Ua��A�I�����V�&�c�ʂ&hJA�L7l��U������([Y��~X:�������?�z}=� nߺ�g�}���sر}>B 04�S/�A��7�ǀ���S�^*`�]C&; �(1Q�7?���Nyvp�ny�/��I%���%|�O�����п���i]8��!��|���L��<R+y��b=l��^Kʆ�� �qc{���X[���� ����{���^���8>����=�2Ξ<��rQ%&'$8��^Edo�t7�oŗ�Q%1�5jq�5�M�b�ʕ�NG�P��8����8n�:a��ML�<�6_^��h�y\�}������ri��&}M�)���h�yT-����b;-���r��?�����?��o���:�930�ӝ���Qn��	^�ӡ���ר���p��������dik�ՕR��W�A�������E��n{�M�Z!�T�yߎa�Zf�EHRr�!��X"+N�+�м|N�h"�С�i8�k�c��`�>�tTw�g�\.��Z''���%M_pn�W[
�]�$��)H������A��7ֽ;���C�GOrJ���^@�̋c�$<�F�j_KEL�J�
"�]��dR�ɚuT�^-Wt]���M��Z��oJ������)_��2	lAH>Vgy�n�h�)_��������U
���`*����������z�Lxlq�z����ڪ�N>��(j�3⢱�&�5�{7���F��$��d��Ci��3�0;y�ңL���$��ؐ�K�v:�y ��"�wQyA�X���Yr��L�!�f���(��������K�`��=(4:8~�
Jr���AT��d��e���y�Id��rY�&���۪�����qĪGD�u�}��oc%��:QIN�ݕ	&g�A<	r�s��:��8��-mK𑆭��oJ��S�t���򹌖�s8��Uܸ~���/`����p��1`��Ko�)q�;{�gO�<��k1��=����~�z�Wʏ:���q��3GpAH v�ͦ���-|�/��;�u�9��ҙ�B땍���Tp;��@���t��ߊ���/���#����[7a��C��H� 50�Ʌe<{�
|�Sx쩧�X�'�'x��W�Y��s�6������)�׷8�E�F<�д�sI�GyrC�ds�ZmQI$�FN'E9��Ѝ9n~�9�w�	H�0���1*Xܔ|DR����l�l":��Q�F��ӔD�����Ũ�qS�������\/>����+7p��q\9}Z6Z��:-6�dGE*f�����NM�,�Ү�@eҲC�m���)n� K�ֵ�)_�Up�5i�]�j�,�/#�)ǰ�ΡE�X74�P����VmA�(N��V1����V�i���qWF���K�P���5˱���J���*��&$h�u��lP��6�I�c�a^`o�!߷�y�E�z���ƀ\������9�~:C%���v5!��_b_��,}��	��ަ��H��&\u���a��3gݱ�o��Ĝ��N%���H��b!���('>��N��Y�FԹ`&�]=� t�Z�Uʕ�Ⱥo��~�y*�ϔ2�����Ƒ�����~���6e*:�����
�ݘC��'�'����c��k7n@�sh-��gcZ(Od{%���Ϊ��Ea�ٚ�t������B���5k�ԧ>��n��al�&lٱ�/�C��\/�ݭ�pk��3�/(���=.Aw��j�O.;�J���LiG���0�S��u8PG�D�5{=Ҫ�lV9t��gu�h�y*F��%�&m�R�ع&��0�<X���c�R ��)��ޜآ&jL���/�M����������O�C�<�2�ޡ�����ࣸ���y�2F�M`]"@��Y�[�4kN�*M�c1�S�Kr͝�8|[�R6����������ψa��^0��H�M��';6��X6wpaj��+�b��r���P/['`m݈����c��ō[����T�>�1�}�\�t�7��_y]5ч%`ؾe�"���"ʲq�zg��q����6���b���rU<���@��qE d��2i�|u��U�3nX4ґ7�`+�xeȆ�!���WD���� �Lj��Ԯ����cb�YS�:�K�
�`���}��߄_n�K��{���~.;���.a�0u�"f�^������(�ASC�!�� ���Ӷ:u�ZW���+�S7q���!��v+�7-M�r�z{��c�9�BMϔ����`tä�5rh����2�Ь�Q��(�l��n[Eg�M�V	i9~�r�\�G�SE�77d�r֖M�y#,Tg��RW�L�5��'�u�<S�\�=L�#R��ʑk�F#�w.n�4�������rkr�Z�� uf��r̚�n��vWV�S�κjK	|�'k��!�rȇ���uW |A�o��+R:o�:xGӸ)�,��� +d���p]��cà�(��nM�P��]#��4� -����&��)k���C#ȥВ��#Z�H1��c��_�qt��O	Y�d7_o#)��|7؃}�(�?pP���_���v}�7��N`d��J��lV��V��Y*��մ.�9nk�\�M8�U�����_���CCΌ;�4��ϕe���A��9��y��&��!��]p��ql��i��3�-�NH�U�y@X�7Z	aVHl���:Ve��OM�����?�5k���'ޏc��:	{�6ly�\�cM�?�m7
 r���YTn�1�[�=�.?�'w&�8sASHS��؝+6sG9�l*�m4=#�H��vPolϏ�����O_������N2�((��镍��w7�����#�v#�&gq��]�yc�7����·ř;zq���}�0�iq��3s�Ig�tTW�ӆ�����T���Q�&V
�m���@���4I�(��`w]CX"�N���u��T�"s?L�Eu�����u_�6Xϣ2������r��ڑM�{�J��A,/,�k_�K4K5���?`���^;�W$ Z�u�v���.Ȇ��@Y���N
2���fũ��3&=��w���������,�cuۑZ�K��Hʽ��K>�BGd �85Jd�[VH������A��C��efY��{��fi��~��B��ŭU+#V�b�8e���H������	:B"�y���f6۪wOb`�b�m�0��{�>h�A�����F�`ڗ�]�lT۽��$�f[��p�7*u�D
=)M	(�j%:b��3:a�r4�LlfД�e!�čCW]|k��:f�V)�u�o����Y���󴇽ۭ`�
K��Ʋ���+��_ʉ3?��f��oH�#�=�m=ο$�5h�S.c��I�F0 (�2���a�[��eM���2��r��%���iA�ob`O�Ƨq]���.`�{�?��gg1-�w|�N�Ė�q�$�+r.I���OqiA�K�f@x�1�a�.3M��� 	~[ç���:��C�w�mW�5$�jv��V:bȌ���@%v��c�C(>�'  �y�3�d�l����9n�����]+
((t#�2.��^���Cϣ.��}��lݎ�ykGQ_��b��� ���1{�#���`�xR�*�]���)'��{ퟢm�ٗ���>���'�����싟��s\�n�'��ƒ�Ϗn���ҥk�KW����<���x�킮x �-Q��Ez`�����۸��C�v�.M_^=��?ǥ$�'J�1>6�T2�۷�Uư&�&A䡌ئNz�Σb�� [�=�����6���ϓ��i�iӡGh�5b�G�[g?�9�ix:r%ޅL�u�F�FAJ���9ϛ[̇"����m� B�\���x~����C��I��W��sѿ�o���uk�ا/=����}�>\��ߺt	��~m{k�F�)�#�b�������ng��h]��w��պ�)��ʶf�ϵB�TZ��XJ�i34Tf-D�Zqz�Ɉ<��8��tv;BbQ�2���H�hGi��v�I`*#�kTK �& ����+�
[�q�P.���S�Ïp��d��b�l��X�{!-�b_�����q�>�3:�d�5��^�!�E��t�H&�<:�l.����\B��]�F��f,Te=����!��w�{����j�>s�ގ���S{��K)+t����/��b^H��j ��+r`R��ϯex��H�!6ыe��}�3�n�p�"���Oat�\�|��7��ޜ��5~yr(4X�>��ӆ |���>���o���6ݳ#k'��[o %A������=�ܚ�F2�A6ǲ��:'�5��$�#���5�yNj#%B�~�� O���/�d�n �Μ|��)�E�x��vŘ5��ؚ��g�o�LK�)!�މJuܛ,=юȏc)4\h�ű̐"-'�}O*�
����K���	�R���o`���زc����t�8�L��]�>�k�����sؼa#��^?��ĩΎ����|�qt�Yڠ������r�8t�s������D�i=�[��ñT�����m�ÕM���a��{��{7ڙؽ��p��O�Ʀ�p7Q�D�7�^ğ�����k���e#&ԩJ˘��㘃%F�
��U؋Z3�cZ ։�����16:a��W��a+E�UY�`��T���uE?7';77�����ƴ[���zӣ���GΌ�f��h=,�u�,�Pp�FõMm��%DM-�|�miڝ�8�M��J�
>��_������`���8}��=�__Z���rͯ`������W��͂ƐX�*�M��s���"�S�8�pXce��Y!�Y�I3�Q2Y}�E	EW������s �&�i��.l_�cA�0:	Wې�����t|��_�y�$��n7�&ʚ2e8}q�g}~N���P�a�q�RK	�\�����ەt��o@YЖy�d��}�FG���Ef���U��
z2��|�#E��9(��P�OsB�n���w�<�������(}5�.���	AÞk���M�I`F�������;_Ʃ�����Zŕo����oc�G�B�$XAɁ8ө�gqa�u�ټO~�S������S��ޠ��R����3�
�ۋ/���ś'N���u��AX�,�NNb�{���{�������q}������o_�V���������3�<���S�%/:ڷ�0���i�����=-M�zq�,��Cb]�����:��L������XfZ:���8r;�@�H�3�t����Y��|s�ԫ��,Д}��)��_����_��\��{���ѣ�6W��=8qܸp�mB�V��鳲�ә:H��Q���F�+���g��}|�?�	�������?�3)�(�鱜 ���D_߆���v��e�I��U������Ё�h���f�1}� �:����~�l\�r_�˯�̹s:�N�W�|&�C�RCJ�46�f�q�+���&u�M�2�q����_�䢰M��1�Iu�v�jd[�:�J+[���u�U���O���������Ֆ�̪N����NG��Dɒ��'͚�Ħ`I��K/@Br|�7?�5#�شo�}}�~�8<�8^}�(�K�R�W�X�͟I%Iz(zM�g�	OV���T{<���>��A+��H�0:4��GE�4� H����
�3i|3Hű�-r�vס$n��\���g�rF�m������+�32���9O1�W�L�2��5Aȕ&���s=��H'7������@uȨ�W�	L�k��~V؛o+��рw��g��<�������D*��P5J`�2�-�Ne%�@L��y}���}͊q��d���4�f�O��*�2�8� ?\�v�i0�Q������{���ʛT3>��xHk�қ��0�Xv?�a	���W�
����$�t/^�܏_@�c|�F�M����$a�x>�5C9̾tK���q9'5�Zd�>�������_�Jnժ�W�uN��La	�9��?�!���o�-�yke�?{Y��N�$A�����,|�
7��=h���t�(��{�,!��CB���]��f�kL�+ `�v�����'�^��]=�������S���V��,b��|�p�M:<���\�sLʞ�eS��Q�뫖q�0�������_�mLȳpSY�y��8v��el�y?.J |��E�l���WE��,
˅�cCÿ!���ר�.1k1����~����~G8�u�eg{$j���{b�}��f��+�`P���,�܅�����+�\m�D���޻�LR��&.O^÷��m\�rY��Z�n\��EoԵՇ���&�6�W��dUs���yZ�~e�MV��@���u.��f�f��)�'b�ө��{���lcS�/FF7'Ѝ�M=n�]�CT���aۗm�7���a%�����X���`�P(`͆u��2���r�y|�S�FV���Q/V� τ}��K�蔫�&X����s��pY����0��Vt�5�l�+��J�3���WG�q����߫ �`y�vM�;$�E����tn脔V1�m��}���0;�t�ǘ�P�03���c�������K#-�]��-5��cH�{�;�{��b$�X%��J��Ze`�~A���Όwu43��>���]���!29�i���ïQ-�4��@���&S$�SY���'�tJ֜�1�4�+Τ���:B�.k)��q���R�ζ���6�V�������+%T5;�AU,��0-�����xZ��/��|#�	�θ5��1#QCr�2��w	fy����F��%l$=v� �?�I%�}�CM�ęg~
?���|`KlE�Lsi��<��cp���7����܋э��\����<�M;��-����	�� $A����࠙l:�B0t7Z���xBy+m� �Hq4���:��U�%Ϥ��v��̛��U��K8ۼ��S��!��C�� \Y�!�W����p�O؎�A���G�B�7$:����:�L�����o�y�:hi�ьD��*�!��ı#�f���,6m�9��m;1y�"��6��� ��}T��`t�]�
n�
���������E��J	�\��ߏ?�������?ǝ�#:S�ɬ8�\��Z�_���}��-K��ڍ�W�N"�9֯�ځ���`��#�4U��0�n\�yL,��e��K8w��f�ڋK8�P�cq"�D�yۆ��	�]��t��Α����iz���dXӺ�D�$�i�W����6���7ً`
t����6�;��Q�Ѷ�@k�f�s\�|0�Vx/��v̹���@3�L�S5N�l���񄶫q��N<��M��{-"h��%��JU�罔s}���O��o�q۹s�$�����Gp���А�^c9+�<GDm���tI�t���</'������&���{�q��ppDkЩc$A��L�C� �ۼ�Tڐ҂&F�rߖ�H3hQ��`Z�F�+q��٨9-A�>H<��Y��X
m�osUqɬ�r�ȓ�s�-��ߛ��D<'�h���:=��̗0�1��#�\��`��-�{80(�V�C��@��?��H�N�ĂvH�㘖�(ȹ�}k�)�$�J������b�y��P�YqZ}��J���)���[s�đܽ�<[Χ��L/l	��ѳ'g�ڈ����ByNuyN��4��.��Y�;mӗ���]r$Mf��e���� _�&�눷c��r����m�7i3�Os����򩌶C���'{�Snʹ1�k�Puy_A�D%�t��~��aӾ~�K?,_-ߜE������hI�նXj���������T����v1-��.ױY�n߮�x�՗����;6_���}�021�� ?�����o�7�Yךy���6N�O�Q�K�7v����������uUL�TE$fV��|ڞ�2�-3��N�A�eFB�d����ub�����vK~W%���R\�1Z��g�T+�f����v�v��u*F�h�I��&(ϝ�̂Œa�k8o]A��%
q� I~N����N���-;}����<>��4FǑ�5�n�v�ܸ�\"��{߃˲>��2�7#�\@mqi4U����$�7����F��//�Z˥S�S^������w�����C")x���M��?�'�^?�1��z�u���^�7����1Kcq~	c���Z׫�+����/��Z���S�fDLڷ#��
{9e'c�d�1:p"C/�n�7�oAME�r��g��� $�`Z�}��u\*y�y�Ӂ�W��7��Tm�P���R�6��(k�H6��n!�*<gqTd�2�gz�(��t�8�8�6Vf{��p�I��5ܦ��5@�G/l��^o"#�h��*F=�7������>�h9l4��G����͘b_fY6(���G4�XIE.�8/�����sy��;$P��II�#�^�v3ӓX�K��WZ3�J��P��h�G��=O ��$��J��^G�/!S[dp��Hۍa��r�qz���.!'ǎ�5C.��� מ�o�k6��K0���W0㖱8uY��J�����p�1������ N��Q�=Y��z	t%Px��?G�R���|��F��u��DA��Z�YD������{e��Q<u�V�����̜4�.�3Jl݊��}(�\���:�[zG�o�Q�o+��4�D,=*����7�l�J:���@!���g���ɣ�mpĘ6N�EBց_�{���4(���ݔ��Lv�@(���D1����/�`+�Z�8�@��
�����Z_g:��!f���d���y(S��%�t��Y|�-[����&�D�$?���`�Cy�����r
��Dl�8��J>�dM%$x̩�����yY�s����������đ�H���\y�[�ډl>�u���#����̨P-˽���>x�)�p��N\��O�&'��;+��h�&��f�I�m7�#B'�#Z$�s��8��u��NWli�>I�$�1�G�F3��m�Fw�;�$�P^V��}#K�r��ґ����v�0���x� ��ZC���
�ʃ1ꉱD*L�˱�&2@s-	p�OB�}��7@����}��~��=X�mf.2��}r �����:��9�]�uj����;N"1���+^��������|���g���~���|��R�S�S'����G��6���1k��y�84�Il��:�k��1AI,�/ �����u��)����X��EZ�bC>� ��L-��i,��{8-MyE�PHT�L�����}e��t#Rd��]J��d�D�11T)�u�a�JMѦ��'�	�c��-@Eb䬲��6[�|4����jT��ה$�1��a
ܜ:pL�9j$4*J�XC@#s������`���m3��N	ǌ�|Nia����ę�T;����ֹ��? ����bR^��r�oKbl�zϡ͞l1^��uk��ӟ�56�-���a���Ѭ�1$A�z$9���jb��n�ܷ��}
VB���AM�_�f^}��ytS�8S���}N�<�(�j��~���װt�
R^V<�t�A��]X��߄�n��!#�H0}�Q�z�>`��r���T]���Z��ă�ۿA��k���a���{���QCm����q��a;qk<�8�jKJ(����d�H?�2�����C��я�����:��s-�(�}����"�a��E��"]�`S/*�ҽ=X3>��05*��{rx��u��Z	�k8�����*���K#����y�m����������:Jrֶ���ɛ��O���J���:���y�>�~?��	P�1�+`
"�=��r�F��9̝��ҕ�����1�tBN�K�`�
��|�i8 $�G!����N�9�+�� ���f%��]��!q�y;�٪��͢��۵
nu��3)A��T�8���RI�'+u�ֻ$��a����i�����|�Y,K�@�d`Cn����i;꘹�ge��y�d4�B�u��s�{C*�V��ӏ�foZ�����)�����)�����ۘ�m3z\��dq	`�ǩj�d]վQ����XקC��gĎ�k�g4e��fj�I����v:��YvzP�k�$�AP��2�SG�u������
U%��2r�k&&p��i�]7��u�P�}c[��_,�t}6SX\~���i9�W$�/��J�F_��/����+�U~�J;t�t���4�r�N����c~��}�E��Q$b讻�����5���"�܊%1$_�Lߞ����]��UH�3����n�GX����X�ţ��M.��g�a��b����F���tLY�*$���w��z�zd�'YFkU�w�)51erSd"C��Z:ϧ,H���qJ�T���*oH�n�}�l$a�j��M���1M���o;�?�C����à֚���M]SJ�[F��M��ی�~	���t�<q��ob`��9��Q���q�q�.[|)���ss�č8�D�e������-ϴ�z#�D�S����'�L�T�駑�y�g?#�W�B��\�M���y�SdЎ˱Ҷ�'��c��!fi�<1ڂn�1��^�V1V�,\qzC�.a��z}9�����6}����#(V @��qv������}e
I/tF~e1nSK%8�����1<� �5�B���xprIUqFz�7Ѓ�=;p���់���`�^��h���f�i;H�=�=�:/��jmI�� ���o��o�=�ݾɻ��Y��C�9v��o�@1�zQei��4ս,�{Hg�8n��%��$�lQ
]��jj�Ր=�߇`�Z�}޶����s�}���&�R��ܟ���5���P5kj�"=	h��{?�r.S�kZ*��f�!�B���F��c��pS�wsZ��8�Y�����������[���<�	V�L�6U0�#�3 �_T�+�K�Z��BB�rU֯ϲg�e���XK�<�kBzl-^?��� �֯߄�������i���p��%�&tN�џ�&�i�:������]m!��p���.N5��^��L���M�A��*�:C"b\�JR���'�]�,�Kr:l�ţ�v,%���l�y5rtq��+���c�,�%h�M�M�"W���eZD]�b�dܰ�3��k��d��Î�ݞ_TY�Q?��~�<��SZ*�}��;�{�c��U|kd�V�nHv�W�K�d����,̎WXBL�j�P���u����}Q�����e�Z��T��kF�O?���^�A�QP⠠E�"��G��Rg1�v�:(a�����\�tY[��� )�A������A��t�֍�Y\M{ak�+��ѩ�"�\+�G�+�U���*?�G�$(�s���8C��3͇��٫DՌ�y.��L�'#Ʃ���B�d�\F�J9��-�CZAMί.hVu��\�
�:��d�!4f�f_������Wڐ�:oK���^X^B�8ݼ��{w��œ'p���o~�K�ЈS�}����r&�O*��섎 �Q5\�;mMM&�>��ǩX��f�J��d����Ǳt�6��^�@J��<Ϣ �z� �?�~ķmC���SԮo��>m1z��V�����w\���oaxσ��t�LL�i���Q8vA�m[��3;w �m'|��z�m�^��koǴ��}c��$�HcQ{Q����F�<(�$IgUu��!���B!L���0��>�yL��}�'��bH��L��ɿϞ�����GQwR�7��)\D2U	����&�% JoZ���;q��1��@'e]�K#)�[���nل�=h	���r]y q+���b�M��F�y"�9Y��]�%@� +�G"���,���H���"Z��ø,no��e-�����k��*>n=�:�/��a�7��J��)G��O<��}wc�}a��%$�{\�?�5=M�X�I�J����������4�WWԹ�y4gn #�M���O4-ArC�dO��\�"��z0%�r`�:x�Cx�װN֬�� H��l\��)���ʕ+a߄�$U��tf�NCO��Q��Q������Y��Ye(=,��7��q�s5�4#�����|%�Q��F��f2�7k )(���b9�"C0A����\�I�mT�
9n�TBC��N`t/t�+�1�7C���6� J��>Q�lB�Z�6�9C�U��M�1�b��-�I�<Ƴ��;lZ7��[�����ĸ��*
�NGw�Ƽ�m�����Դ��}�N�3���wZS�|�.���W��+���w��ī���=��ǼV-y��o� ���EB<G��L�uV��L�J�K'N���^�)�	J�'�u�h���R'�#U&.p.L�ԯbQ/0�c�7�6k[��)�Ú�8�~2��s�	"�<a'���M�|+7d�D���ݘ��Kf���b����ϊ�Ɉ3�������[��IM���47O���Z��F�Q�5m�u�Uͱ���&
7jr�ʹ���`�^���b���~{ �✖�Y���������䞤�+H�-�杻qdqiA��FSդ������y�r��ړ�*�5�Šdbh�9����v6=:��Sߔ�� �(Ȫ�����=�,��b��h���W�f�&bd����A��Qz�,z>���������~���8� �8;ӏ�.�/�Wo���1�O^��(�˳�w����З�=��S��h��1H�8��!��&��?��nq��x���s��1��c�������a@I�=���ߚƚB�\R7�Y���I!ʹ
:��mo�hp �������Hem-ˣL�?�7Ku�	�H��t��:�����8�n/�)9�Ag�JcA�㚝;!��%q���Ez�����1��n+@:�*��N��v�m]��,�]d�h��О�"�Y�[gY�� ʔ��R���`W0��>��/����X�����dM��b�&4�|�
쓯!c	�#�쒭�z-��p��li55��q�qQ��"p _\��>���b�D��������7�n�rS8����_�ˇ�<rZ�-��+a���[�����P�MIh���%�g�ڥ6��+�W��MB\oo_���MK�E�ڐu��y�A|�1��(Fi��N��L y<,B���9��lWaL|̐`I���=+һ�� ���\o$9ˎ�:�0��-���,9��%ᑟR),���]|᷿���!=�vΟFlb[����6Ȟ).d�z�Za�C=C�?��?cID�)�����?������_�ׯ�C�B��t:cٝ`�?���:���ٵ�[���;���[d��2�Ȇ�H �2���I<��3(��,�-,�ZԴ:I&$����S�)�A��6=���`���22�Y�沠��-+��N[J*zN�&sB�pF�K�H�I��ƺ��{����\����-I@�k�J��	�~[�ءD*�_2AJƀ�-v$�PS�F�l4����Lɥ����V���B#q��y���X�G��l���b8��KZ
 �HR�*���������6ݥR���A��.�=�tK��e�r}ԩvŨ�h(����W'B�$�^��uqi:����-�;+�G{hk�K�������,m�:��iȵ�	BK2#ѩ!�n`\��>t�}��q��=!s�W��9&HH
�zz��,��\�µ�>��[�,���h ;4��~�>�6�Ư�!礣(%�i.,a��p�����8�8��ދ5{�b쑇��@~X��gY���}&�N��n�G�ӬU	N���������zd"���{+.�q�VON_o��>��c�Y{pk�=(?�5&K�[�c7 r%	4��3X#�#mK )^��3N�Q)�Z��y`/�,�F��C�`����ۻ�7.ߖ���� ���A$;KJx���P�8�LZ�A�I9v�+&HU~���Ȉf�4��>5����7��ί��}���{�/h4�� �a��g�d�,/�T�\vGV*���/H%�JŊ,�c�.;�ˑ��"Y҈��g8$A  ��wt��oo_��9��}�*q~�Qn�+�����������9��zɉ
�����o�%?����H5i�b�u��57QJu06�����w���42�*���5�O8:`��,13U��ǌ��¡�^ǡ�/�����_Deb��1��Н,<x�o��6����m�0�J'̹�2��ŕ"Թ9i�gIc��,�6�l
0&� �k����󤒺Ξ�F&�g�,�=�F�$�C?��a��G����,�I�
�+w\o4����mY���@��lb�v�X횎�H� �[����hT-"�s��9�}m�[f32X�6B�*���Q��R�k����&.|o���m�%F�>2�5�Se|��9�]πs��|���J0K�'31H�OFwg���~�W	����f/��t���W��mTѓ&}/ų��О�/[[�;�O�-U�F�_.��>���%"P�DSذ��O/^�7�,=�TщX��SA����M_�,�-U2�J�R��J�P�8� 9��b1gD#*Oi�D�me�.��.ml����m��yx��b*XB��g�D�/��.�L�W�_�F)W@��G#����������*���6d�e���j3����x z����J��뭞!v]4�Y��ct�!j46�v�6��wx�^\�t��������6O�Cqe���t�-~f���0ؐ�l�I��C�ƥVopmilh�Q:|}�=���U)uxG~���%:5�����:��?m�XH���zwm7��N������xabF��e0���K�~#?��K)�&�&F��K�#�k��"�͠�)lְ���_Z@QN��닎�F=3<���¼I��-�����ч��5<��LÿÀg���?��ɟ��H�9a��^�J'�"��~�����4,���y6�w�;y��f.���&fR΋�fQz�E�GF�Yc�w�:p�$J{`��o�G�.�P��1C	�t�����%�\koa��
�^d41�*1}��&3�_*c̮�̾��>{	�_Cy�_Cur
O�lk�u��5ҘW�2��^ϥ�|v�!g��)p��؁� ]�9�`N}����6:O����^�61�����=_hf�-FiM�]f������C���i\	�K:p��UZ͒/1 i�&��sӓ�8�կᇟ^1��8_��Q���Zk�k���w��5�>���f�k-{F6�3�9r�I����:���3�>�� h���M��hfub,}ӭ��VALߨV=�e�0�\֪�z͂u��o�S�ۤ�t��9�=޾{��v�u�����v=D$�����k�Eʍ���C�:���EX�~�h��Fz����GA;_m��R���Vi�$ݫq���}:�	:��qTFư�����G[~�׷P�=��w����卍ײc�7x]�K����H0HU��Y�z&z�f8�P�0��H�L"1y���b��eqCt(�=��A0:�� �L>c�ԉ��?�ͨ����
�2�N���7�Rթ�9`
��Ы�@#r���;u��������R.�Z)�A0�IS�W�YY���k2��F늘���9Z!؍��&���3s.�n�mNY\���Ms�3��4ŤV!�&�QH笿��ء�@#�7��(
v��H�+�deD���ő�	m��$�LX�p��Z�`��;\)1��S�p��0��n��eu�	���G�F(��n.?1��{��{Ү���Ƥ��@��v%Ke��t�5�܃ԋ���Z���/�_��h9!�xUy���.!���#��Fp�$D��{����? ���=G���nf�a���Z{��}���<��Yưʾ	�w��S�e ���P����
��ѷ��q�9�*'m�:�Z�h"�&��+W�:1�������x����W���Ϯ�ŀ1���gѣC_}�
�Gj���H��+�ut��C�6��G�"�`b����R~u�Ն��6y����+l=^���?�q:�R�G���,���dΖZ�1�����5<��	b���!d ������X{�d���{3Eg�7��Ud���<���u<?_���k�x���Vǧ?��x��
�ێO�a�k�a� �'l���e�
SH&���=�`����[,>{�^�Z��f�{�T@ˌuG�<�ӣ�������L;f�>���4�Ç�q��9�0�;�:�R�S�LD=��cw̎	ҕ���@�α�Ō�*�J�00i�\.9Q&|O�h��.���/.;��gk7���LN�V���!�,G��(!Q �G�L ;���D�Q��@�Xlh���GL�������0z�3�;�����V�(�J�q}��U�Hq=����m#E��@w|�.�{զj��
�:��
���E�6�,}��٣�Z��2	�\���CiF��g��K�o�񳗥?�]#�3�t"��;�l�pl�Iv��'H� f����k��z"O��M�b�,�����>���*�4��?�ȖE��#(���[q��_�t�0Q(J��"�rN"���U�#�ba�R��q�����C��ͫ�\�@-*��Tʍ'��D�""��H]�ҩ��qVVgt����f����&i��J̙:7���O��y�'�x. ��JCҌ=7�. ����鞌�F1�DD��T��{8�ML�R�Y@�0�czj޼��~�}����U��M �љ݆e�ܳ;k�>h`Zj�����I��Y�D�v� <YB$%22�8/�q�?n%��İ�0��拸C�X�Km���/F�dOβ���ڃ�h^�����s3Q$�x�2������{�6`*��Bf]���q�p�i�k�Bi4[w�}�*����\E��̋�F���w
���̝� ��N"���з	�6��h����O�?�cvە7(�A&G1z� �w��������-욵�^��I/�c��%�~�Ʀwcױ�>���??��W����(���~�%x/���̦�6c@�K��k7�,3��͛��L$�l]�C����8�*=�<��)��9��ưb�Y�n�N�J;���|�6_��CZMe��+b��if̳�-��@ �t|7s�K��Y�45ˠ��r�d{���;���=g�>���qMcY|�M�{���mўd'�q�K_��;�P���V1��k���,�����~K�M�4
��Y:J:�����v�F�����#q������U1���[�Hs��jjG%���z�시bܝѝz���l�@�!!��W%�*4ڵFv�\[��}�1<4d5˺��;l�1	�ed�C�t׍C��9{Q1��6�j���E�L7fDI����{]f�.q>I����k8�0[��xm�Af]m+�Y�̠����}X�{��/_�i<_���·�^��0��3ɥ��,��s����~٩��K�"��dJ�#�7.'}:���,erY���axt�rƹl&
*��Ʌ��y:�D��@ �V�͝�}��y��W.�9s��,RY�s�]��r���	k�K��S�s3���Am���q�5~��t��dU6K�/a=���@���X�t�A�"��p�vL(����kt�tJ:(5)Nif��u�Ut�f_�Tlmmc}}� A*K���z�2R�)Ĭ�'.O�o�,;"U 6Pe�*�f�S����{�\1����,,�arr�9���(J4�
	
�C����`��fĄrW`��%=��g�I�����:<t�h/�͠�I�n��b��9f�]^�ީ�V�U`$�	��<�*׻Q��)�q
������A�W��,H��h�o��x���?��a�C�7-��)�Jш���%k8�~��:��*�(�ZR��Y�W\}�0�� ��:�Ⱦ�oWv�gk����]������n&���;���-Xou+d?�	!}�0�@/�SY~���J��0y�(6`$�4��,�{f�P;hݼ�q>�d�1Jcs���	r�KeT��*���4���p�n���.b��3(�ۅ�ѾpՄwb��֫�v4���uR�*V�%$j��ȱp_n�9vf&��Ͻ��石����G�޺��~��z�2�׬ɟ��K��x��|�M`�,R]U��9~��O�뵱��s�t�����p۵��b|�5���{�/0s�9r�0�gf�XG\�*ϝ��?|�[ĸ��?�H;�Ѯs��Vs�Zu�� JY-�z*����
�t��.L� �ݨ�.�\U�tj^�ox19J�G�3:���Ա��w�����L^,B�;��Vp� ^�?b��̳~G `D��{�S��U#x�=��v����>?����d��'�����f�q�u�IQ����V��u� 3{g�Ȋy�@������a�&�y�k=pK�ny���D�|5�{���j�3�Գ���9t+m{n��[��Ȧ^�����O���4�,,O�B;_F_%hn�N��b9i�Ԓ�Tv~��asmŐ蝦o�//t|��+�S1[�[OY+!��,�zܞq\X����<��	���@A���c�F��nI��;hvz��H��O#M'�g�R�T\�?�W}n�a�\$F�q2:�흺�ʍP"�l�<���l4Z�I� �t��	D����W�<4U;�
HtX�x��zF����E<e-���(cn[A�m�w:������������*ν�~���"� �4���޽Fj!�-:���6�e�M�Y93��� ]�Fr��S^�/}�)F�"��\�3;k���z&""څﾃ��{q`z��󢄵��H=M�-Z�DO���p�F��r�6�?���=F#���h(��b�w��c�Џ�(���i�9�9�d�m�H�̑mloo�F�_�$og�X�v���))�1{�0@�""�>�W�=&��A��"Zg�b��1:���"��?4��ݻQf���e�7�Iv��Z��c-z��P��.r\�:���ְHg�U�TA�*R�	՘r,�M��]�H�xa�����H�}�44���2�>~%�����Ѯ:���o�^`�0:T>3�co~��4��,-a��u�0��k�NO���߼��1�m �l4��>�#6wC�5�'�����2�{Ӎ�psJ���9l?x���E���G���h�D����^Ǎ��QE�I����=P ����O��V���r���gJj�v��,�H���y'{���"c�S�y�GR��p�ʦ�lb��@��S��C�N����{E��lXf�7vX�\B*"��"@��>hZ29S��ȧ=���z�@l��6ǂ]#�w�+�_�D�验��.��s��z�
����F�DKb�ԁI�t�[D�k�i����v��s}�W^{�����>�m����n��-c��1,ߛC�qkck�La��\��[��������������??[��gΡ#"M�7������'s��GSƗ/�8>�V���� �M�E�r^W�|��7���$#�����-$��'�&`E٩ƨ$��;Y�{QF�P��,m�(�b�t�bn��Q��Ļ=G�(%�f[�;�_Ɵ�&��W5*�6f�kd%��@�P�j�b�LQ�v������Ƕ������E��޼�rp���ul�Gy��Nr�E��PŜ�f���2 \��K�VsLRL���U���)��+��NV��k�ű�d��?�c<�����(N;U>��n<�y=��D.��f�J���J�A���ߢs�|�������2K1j5���?�֮\é�']����1WQQ˂�2��̨�@c�J*�k�9'Q�Ű~�ʷ�"��Ge))�v���>�����x]q��U�0R�6
�T��]����9�i[��q��>���{#F�9����E����s����%F�fw�w�A�W�`O��H�P98�ՇW0~hJG� d@�r�.��NR�����F�?�=���`�%f�����7����>��{*nE��64�~`/��!(}���k��F�fϿ��ĝ�b��������iEq<z��%x�±�l��O��:
����n�$Jc<��sX�p	��Ex�2&}8@\/ck�'�.���epA/�G?xK|q�oB�'M�#�,�0R
�[�y&�-Hu�\��F{_z��Q�o?�ޙ�(j�N���c}����gv�`7��И�F�t&���X���y�]w�����Uo����l7��6B)������{�	�(%,�ﻜ��{����L�8 �s�.+OD൮Sĉ9�6�|M��m�9�F+K�)s���T�G�bZ��>g���L�Y����'�/p������6y0Ҧv$�SY_�C64j%(�H[�aex���]>ϝ�o�g|��I�*U��6l��m1F�T��F�z������ݯ�\���Gzz������;�v��붊^�+l޾K�UZM�8�}:3t�|�8�����>5�q���xcgې�/��9@H��Vu�U�SnX��2�7�/��iw���n��!D�b�qܼ���-:BT)�e�E�ؘ��d��Qr�*��)�����H�07�}��^��CG������<�[�����{��U	M��,#k��W�����!p(�
̦���w���/�A�?��b;2B*�
$�e&�V\|ަ��2�~�զ�1�JY�$Ƹ� �)X�B��|!��L{�GPߪa��*��S	0��F��+��׮���*J<�Z11k��ٓhK��i����}\}�[8�lt��q�o&J#"���+��~�Τ���Z4'��"Z/>6\%�U9���z��i�'��>|0��s�`��I��w�X���ڭ[�7V�;>��瞩�0P�L{ת���R��{ �kS�����X��!�������O�48�%Ts�d����阸��c}�	=�?�V�m0��֕�o4��ُ}�}��/�8:�����;X����#���V���V��������w��S��Nw����9�*���	����(4�����;u>��:�ܺ�9<ȡ��g��sU�:<�]�|�{�mz!#0�*M�������iX�sk�."׭sM�ơ�>t �W^�:3����_Ʊ8���*�*
r�1�Գ��,ܽ��71!I^:�<����3HJ8!�C/��&��
�d�A����@�~�5�޸�Q�3cc�䦊m�\��3�?���`��)�I��p08rc���y��l\�r�)XI��h��d�N;'yQcZ�����#R�n�U�%��㤐�%lVc�Y7�b̕�����UP;O2�<�"�]PO�A�^I��T��[،^�a�c�R� _A�ڍ�Om�Nv(]�X ߏ�ۍDg ���i�ʡ�z�g�X�7�kcH�+������!������Ҷ`�q��%\|�3�����~t�;M����8V��P9| O�\E��/���ד��[�~w��bEL$�}={݋�Y2>�Z����i�-�~K����GX�,n�(n��H4rS޾v�[湶�f��q<(;����-]F��wT�6%�u�@yv���I�sE���	Ѥ�x��a}dTPd�i7-�TK6��/�b�A�9ӚE�5f�͖C������y̮͡�0�P�����<�Y��1T-B�	7�z�i�:3�$�P��:�6����8J�a<ij�g��]gv�g4N�>4��r���1)���ܹP�Fo�i�2�4� H�b�b_󦦝�ޟ ���d���$.^����Ǒ��L��������F}my~~}y��i���ݠa��TY5�SGeeՅE̽�MF�d���5�k���w�}���IC���KW�l*Y'�:�7��ff�w��t�Yi�7ih���^��U��4U������ъ*�6�R��r��J����.a��_�c��U~�'��K[�{���:
��s�<�a[,�p��t�S�p��;�������{��N���5�s�O�tZ�P��"��}�f&3z�����]����n S�a���*�i��3w�]�HO@orAqĪ ?�!��7�i�@�Py��4���P�+�`ql�^�į��%�Ʉ����Z��^:�G��r6j�Lz6ff�*F��ǣK�����8��c�gf���ؙ��NNctb
/�y;O���Nŏg�X7���KYN�u|�"��D	(�MXGS�����>_�~^�@�)�����BG����9�;v#���p�N�y��s���w�XЍ۷p��sN*I+���	�C:��浵:��c���HU4���� e���I������Mh6�`d��鴑EY�,����HX�75[��]"aL�Ɲ.a&���7���`W`�v�e6L�7�/�K�6���Z�mj�5�M��U�'=T�~��@[��@�Ѳ
d&�ut�;5���i�2"��9(SL�=�YtI�
 �{��ł(��Z=:{Z;O
���~�]/^ŉ�_�=WlJa���rs��:�mXwb�	��5?�O�-?��Y3��*h�,����o�K���Y�z�:l$A�|譀[a�����ۅ��f��ᰨ�bB�TRB�f���
v�w�9̈́+��3�u�C�+��ge-�s��W%��so;$��{�9ommX���y�ה3����2rn�B��6���V$��h3̌U��F�ss�H��ŋ�\���d|x�2}1@�1�{O����jca*q�i�
4��μ]����Tbuy	wo�`�޵J�J�#c�\�e�#r�F�*#��1�a��k-Ĝ����g������yϓ�e��|�^�z/�W� *e�󐱷-޼�:�ۋ+��B���C�nE8�)O�&h�?��;���Y��������֯V����vM�e�nh�#ɔg5���8�D1�ָ�ډ�9�F�t��%�.@��,����z����y���K.2��u{/�u��ѿ�Ǭ}��'h��1�Bt�x� ��&�N��P�\��0ssh޽����^�7��@�*eYl]����o"dp4��	�?f�KX�Ǝָ�����DesE�N&�ï������*�$�S?_����~���m�}��>���0��M$7wL�El_��N�T�V�T����U���	���F���jWc�q�0@3t#OL�����0��J�;���,��>���O`��q�8�	V��\Ho�_����T�6ۑD�1G��$�p%`ߡW�x��MY�.�Viˇ��C_8�-:�4�43��N5��}�����[�+�G�mq� "O�M&t"ĸ�v������SI�T�&g�s/<���F��<��J%s��{d������x6/�݌��TA0e7�D��G��{�����?��7�c����|?a^�}��5�ފ�}ʤ�8t�a�T_[^�qD�h뗫)ڮm�'׬3�L�C�gϘژ�MXbX���XSG�O��[Mt=f�t�������wp��AN�Z����3��m<Fqt͇�Ue($�8�u��{��Ɛ���J?K_ϤCO�@o�|o�9��՘���1�g��7�h��Cnҡ1Crf�癙뀪��>'o-�����ۀ�8!@u&D�`��*qu�Vr�]B
�֮mR�������FFG�z5��r]�Z��Ȉ9�<�@Fэ���t�H%�<��X]^^6���	��w���D�m�k?��)�=^�E:M��i�Ejg�[�v=�LЈ�0����S�y/t��qK�--�F~�� S������Ub�h\�ODs����N2��	�� ��������a���\��"N�y��^Ƨ�H����4�Z�9�k;�g���-#��Ml=y���$�����}��m����/c��_�8�N�@f9R���d��xS"b�9��@�p�l����WW#i~߀\^���%)�i���5�!&7f�yiүn�ѻg1;{1̓���à��I�An��aZZC�F۫�=�����ѭ���:��e����WQl�ȴzVR/���3�^1Lb��
:\���0|�9~L�_ǝ}��N�
�����.桵�,-S®�y�1��|�ҹ�h�z</~��Xˍ%���nSf�(�6���������j�o�,�p������l곻0��W�av=��k�~�*�$J1�	$�[�kX�zqO��$B8�r	�����y�!�g�������8S�@ ���ڷA�i*H�M��"��{ۋ�R5���_��j����3�%�����.�:�W<�$W����.z&G���x�苘��@51aS-���գ6�d8퇸�B{��w�X"�����k\5�@Y�TA�Q� 5��&�
��}���aF��)+۠������h��LV���ٵV�g�1k����E��K�/*�Mu�����ܾq�t :|v���� �\�Q�ҽ�#J�R�#��{�i�ߔ��m��g;Қ�UD?��HՊ���g`{��qc׳`��'��\��m��6o>��R7���'R�����n�3��ϖ`�3���o��s��5��v����j��ӳM�`vp���q; ^�n����Ĺ?d�;g����8�b�Dɚ���H�R�X�P���E�"O�LE�;�+�
��㵨O�C�����9�9٦V?L�x�H8R6��֟�(�����=t]r�gΜ�����G?z7n^�'���|��M���o�����)~�Ko��_�*�?x�yf:���on`�©�N��7^ǥ���L���;�A���r�l��31+�������:�B�[$�9I� ��MO@?�S�4���0�2s[a)ū�X[�\Ø�އqo�0�w�_�jZ��R�� ;���Q4����Lsy�h V��Q�,�Ъ�dޡ�\<0Z����q�t�߸�M��g����sN��rÄ�"9��[w����{ѐ�	�0��s�c���X�O`�/�%:uf���{t
�if�̈Cf�B����Ŏ���7:g"���#<��Y�2��D7f�cu�Ur����\_]���0y� ��ڇ@���
�;8�f&���b��`�E�����f���Q�;Kg�ݸ�ץ^��Ј��yJ�l�{�p|72�#�-�{�*2��b�AQ�c�������n�:H��k���?j;t�R�=H�M��^���pm�
b��^=��5�˟[�4����O�έ�X;{y�]��B�5HLD�*�iJƬ\�.簘�-��T����������F��(SD9r���f�;(q�%�9cų��o{���{w1�k�*Q;F��3W�? ]2vcJY����)+*�U+�d�E�*����G�Z-Y�a������-E�i�X����KW}�(��{z��L�i�U�TaLD���8f���,�q�j���z�|n�|ݠ���c�2��rŦi=f�ǵO����Dl�	Cч�{��k��
|gD:�b��/��ɉ˶� @�N`�H��^kcgs�F&�\���/��]&��5V���ٸa���kd���VV�z�?;�I����4���E�����_B�F�y�5�q$��N�F+t�t �|������0����)P��05j����~���*�t�4�����t�Dl�H��RV6�!h��}��$�_ʦՏ2Q���}YV�>�����{{�t��4�������+羰�h��/~���O.���Ǖ�>�_������#���[x���]�����at|�ԡT.;t�0v��M��sϟF�ZƕO>1�%f�B�J�MJ�RHM��[L����TC9��#��WE�	�D�T2)������z�2^���}7��g�*�P(�:6��#8`0�
"�y�0��>w�V��������t���T
�$bt�i^W��o�
a����<�	��^$+gF]��d���^i��t�a�zQ���%t��J���e�5Qv� �*�3�m:d�?[�ڗ��;%t�E�Y�dZ�}�d�ό8�u�uC�?x�Op�O�=�j���$7$�3Cץ#�yd:���M:��o��қ�Q��C��@Hgx$[�LصgQ�g�P�\���nc�019n��76��#֫�>C߽��<���N�0��{g������Ve���l����@Vm��l��1:��Ait�^}�o}ς�����$E<$�V�Crk�+$}�@	��i~v�[���O�?s�WO��O|sW����F�p�1
����kD�7<��AK|]�+�w7P[[E��{2��F��-�g���*f0u� nݿ�YZR�K�����5U����i/��Ҳ��ꥫ�g��� ȍY 3���%���#N�h<��[2�h�m|,��,�c�4���Zp�6�����WY�;���sI�km5�酪e���"���w���nrȱ �$x�+9Q9\g9�vdV#�0x�����^�RB2�6@�6�[��s|z�Ͽ���e#\j[UV��(���z���:��z�vi�]7!��$���+ev��}�k7C���0mKLD?z�i���.���ȍ�a��HI�|a۫A�~���wz���J���5��o�K<_ϔCw��Ff�Ż��K�V����px>S��P�ʬ�X崩j�m��AT���n������Q�ʹ3I��2����LU��BcFr�*C�Kd(rb:���xT�&� cP6W$�*�4�5sZ�m#'���x��p�E��h\���ѣ��Js*�˩��_Fu�����c������g^~?��?�CGO���o�����/��/⥗^�ӿ�7��J����������/�����mX&ݷv�����KD�݈��3e���D%B
��T�P �ʔy�����}�!^���$#��D-�Y��hDԧk����X]A���t}EJ�uxH�=':\���%�)nf���ʰ4�\om(�u ,:���c��H����f����dؘ��Ջev�H�1d��3�]��UQHؘR�f�E���]��%�̚X @���2�YA�P<u^7�ė�������m^�@��-<8�}�������qˈ�S�"
�r�j�6�g��
,�4V��]\��k��Et�<�L"���53����R2���j���*&��Hr���\A���E%��6}mb�l��"ƪU:�!`y;��"�dŮg�m���a	/�W%.��}���?0���4�U�ހ�D���M5���@/yER�_)��s$,:Q�v��Aqb7f����;߆����Jʪ҅FCf~����ЩS\Ϧ����[���"�ղ��c����������MLNh���<�¤I���9C���5�\�3й��1Ź=�DU���J���;qc�3�h舣l��?��e����J^��{z�4���ݻ����^UɫT�F��l�2�Q�҉��׏��WO)M�
�E��bҵ�B�-טl��N�o��A}`�T�R����T�V.�\K2m� N^y������-1Jz�c��XV�3�7�����O��Ԣ�j��a����VƏ�P�Ǳ-���n]���G��!f��� �_>�o/�Anx���N#�h��Ē�f%;��{x���g'K���=�0t�X�?�뵇�,q�%����)㈧ml(t��1޽s[��,��@ "2�8�b둙�a�z��1�}7�f���6��~}�.ꗛ�W�CZ�$��]�Ц]dF�_�3ũ�/zT�%��SQ�r��d��fu؄x�z����[_�/�d�Q����C�U_�qӪ���5��W��u�O���?�g����������k���O�}��'�x�����6�r��a�� n1k�Wtl��O��FMW\``'^���E��	�!�� ��bV-İz��|�2�R)�͍���2��'�G�TE;��n�a�=d;X_Z�ۿ��ȧ�(ӡ���I�
 c��5��d�&�Ynk	�w����]��7�h%����P��\`����Ϲ�o��x���{� Ӗ�>��r������HF�X���?�7��FA^tp}O|����P����)��?;I���n->��KX�}�|�I:��T��}#��1-�j��(�m��%b:T�%��~�R!��ūH�/+�����2�H��|�H;�o��ַ(پt��9d�t���M��׻X��{&��ݸ�2�U\�b�3Axe{���9�l���Z�������!$�V��UK�=�;��3�nn���h���߆���
���ݾ��?�6��SȬ��33Hi\P��~��QZ|�kw�m�]������ZFУj� ��c��9�؏�n�Z�i'�%���8��9�1��~���fV�~��9b���8�ׁ)0��{Kճ��!�^�DG�q!���ёQ��º�M2�N��ptTr~
�M3׌�N�M1+u��$O��҄���]�nz�Uq��{6����h����N9�Ӳ�6Ͻ��f���8��)<�[��B��Se�*��$���!��3��Y{�����G��-炇�j����g@z��>9אA�����D:�w�޶I��5M	�>�sԤt�$�S�Gr��5��j:�����x���xvh`�)��P�7r`K/��ZŔ/3�d���x	ˀ�Gt����۷nبE�we^S2R�9�W���n(�(�0�DD:��H%JI��D!�I�{�!)bi0�m�������v��A��z�V�Sɚ�M�3�ؔ��у��U� ��˘����=h�./�b�����~�wo��&�����;tP��_�k�ݿ�w��3�������a�:��xO/�
�_���K��=t
��QX�?|�4G����4��xhi��js�����_�ߑ�J�sVUih������o7�ϭ�����(�9ޏ�2��W.��^�z�Y�v��-���FC۷,}��7�Q:�>�����1�yRiFA#h4�%|;��?6^vS뒦9_�C�V�f׹G�����d�4��k"�kbt�j� -��{��uo2�ڛi�̺*�:;[H���]����c��W"�uUf�\K#fY���g�)����Q����*:��(L$QCo����(��6���o���U��<ت�y��&B�n�!�ա�����{t���K�H�(Fg ��y�~�i����;غp���
�j��%4����2��.����e�a�4�h4ϦA�P�����.����ָ�J��P��4���b�ϲ��A���!6��l���lTN=����}��}d )l��F'&��c�0����s�Q{6aѵ�\�u?����J��i���s�[��L����������)���t㡓;5���X�!�d�U�t6�ĤQKc߾��ٵ�0?�{�K�LyMΨD�@X�_oE��S
Xϲy��d
Y�����g����¼),�*��� v�=�L��{`����GP�C�䰭Ӷ�iӒt�ci<�w�>�����1I*{��}��u
s�������h>'U)�׶J�������D,t���H7ŠLA$[�S^l+���=!��t_�˯�-X�iԁ���{{��f^�*�]���0SIӳ�d�5��ڪ͞��3��u�]�:%8p�F���ۈ	Sr�p}���b�bQ.jsmloѡ��})�Ű��A��ٌv����_����Z__��>::�Ey��t}m��E.Й���j%i RpK<�v��M�ٔ1�E�y ;��/bss�Z��柘�����_�g�/�－��7��7V��q��^����0���/��o������:z��5����ߵ�<|��{��Jݫ#�hC/�7>|Q�f4�+�K�Yf��������˯�3W5"_�:�6�&�^���ƞQ���̪\��Jp��XꜼ��q�xȳt���f=��m�,�6�0ꠣV��tE0^��p[�H*3.�<q�Tgs�L'-�d&�������z���2� d��x�ku�t4D���
��I$���4��۫�m�J�B��Wب\?蠭�-��A�(�Zbi�
2�`zBs9�K4o"@��j$�f=k�4����f�K:����C3:+�qMJR����ݩoH�М��U��z"�N��@�6:�mw}I����i�Qk���U%� O�A�C��u%`��mS��y�]��� G��M
W!ކ�MjI�T��m�[+q�����Ͼ��->�5rUdU̯�`��Q�+�Cy4���7�7,�z��Z{�iQ ��D���I	+	051m ������F�)Y�&�e@�!Z�b���N1;���ʲ������+8}�Q�>y�dwll9J��������З�Zr�M�$���$���/�99�?+�C�y�Zc��ʷL4Jv�X*Yk�ȑ�g�~\�q+L�t��) 9�������L�k{E:U�iD2��E׋�aZ6&�?��5	gڪ�	��Yu�����Nx��7o�^���?m�L�RAG�	�#i"Qa�Aߑxf��w�W2HB���gơ�����iTvw�^���&+#�4����I}z��u��躕td{}'0 �l�^�h<�c+�ۼ� �
�	���t7�IL`��}V�z<?oQ��rm�={fMRT�O�X*`rr��n��l�33�{瞕�L^U��}�e�4&����k�,�V���:�Q��_��8��@�~+�/���{���I�X\��3��!���O����#��jh7��ȱc8Oc��@H�1��T�Z�)��(����_L�5S���C`�/9:O�(�"J2��#�����'F��1����2�hS���p���ۼޖ!�E��6�־ehA�t�˅�t�����1GX����9��{q�mjF^��s(�,3fo��b)��N2(�����9T}�t�1Wx���R�2��9�]��y�G�de�?aل��xĬ��3�x1l����I�:y��{u7	�]����n��Ȭ8�C�hȳB-3�)��̡̯M��+1��G��icm-����+��8h4�M�xF�k��)���)1(��`��l�z��z��=.��D���a�i(C��w��n�Y����q��N����7���!����`�D�dB%	�P)5��O"=}!�N�X��޹^
<ā�O���}��A��dt�>>��{O�di�B4f)G��~����z���v�
�c������
U�$Q�^�)�h��'�_��,����]�ؤ=(�8����P�8�\�Ui�ߠ�*�*x��8���w�6>�9v��e�"�p��M����9;1�g��4o.�m�νE����f��()�D"m�r!����m�?�E�<24��M)���".|r��0L[���(��cڐk�|��X*��iK{A���$" �Z~I�J|����%"'=��$���F����G,���Wd�<ka<m�h����vJ��#��.�1	��w	�?����_�����_όC7���.�������҅܌�H��<c=.�xön�D]Q���z=�xc��q=+"5��Dr�&1�HT,����ef5)c[z���֬l�n6-2�f����������p"Л�eB�;�Ә���G�{����Yt�ޒq�s��!
��]�Z����n˞��ۏ��؏�����wߵ~������&J�
>x��8r�0f��x8��Sp�;2�S/�DG?��-F������D#ا����r5/. ��2�3�^�k%f��4$)~�A���2ffs6fT�
��<e�͂ 7�I�<eU�9t8�n��o�p��M�4;-{W�q��$(�V2�������ϛ"��3n���m��0�;Wp�7+q��C7~���]����o%�27�.�yd�4f%�ft�|?�O�gY�e�~m�^y� Y�w�cB��p�X����6�_�	�d�=�`���h:���Cr|m��q�׳���->C�x�Bg�%Y��� ��64�g6���9�ϸP�L$���Οg�_��j��;�:3/e���C;��!i<��}:J䕝C���f���Z�÷j���IjB�KX����t┗z^��Ћn��g�A�f�6f�-�:�#����[�.�o1:��(� ڃx*�,�h6&iN��wy��m�9F;�b${*��V\�s&~D&���{ZV�����uV�Z���8�ҋ�^��|���C���O(�����W��R`.�!R���5�Qh�&�ᰁ=��~��MrX�>�f�ΖJ��f�n� �TEu�L[��U�PԬ��l~s}%:sMଭ�Zu����xH�j��[���?s��lq�Uyr�r�b�$Iqߏ�{�ԫ��mJ �#���zn�X��H��Z~���s��V�w�!;|���/͡7����'��*�>�j1�m�6M�6\�q�T���_�4>��Ʃ�<3�!:�|֑>�B�?v m\#4���A�\�l���tl�*�9�yO� �C��w��nF͋���q�I�1�������.]B�R�J�eN���v����*������}{@��é]_���:�:�ڰ��݋��g�4�Y㎞R��T:���;��;1�����8�?��|�-|�z~��I�
������׿��d_d��g��ՕRNAH��@�t��-�aE]�z��D����|?�h8>*�7�9jH�"l��ҡ/af��qL����J�Wʠ�,��
�Ӈ�Ez�0���oh�Y1���/������8�%�19���ΠFó��9��J��CWe+�:5b���C34`y+��f�0Z^{Ϩc��X�r�w
"Ui�3$.0�P:y�f�h�=�buf�5#��ǻh1�*~��H<���u����4�~а9y��5������e��O�n�G��"~��f���4P:�F^}��L���&����(�6i�3r���Mc�����kf��F�ｸ��*�4�%�����9U$L!�s�Q޿��u_cO60DgI\�=6��MA�9i�yN2Xk'����|o_��������xf��9����[��h��0p8
�0Q5ɏ�.�CW��4���%��mjz��n��|e�Y{��dt\��'|�=i��A�uWv����O�HNTe0p�.������s�5Q�Tٮ�zskː�MNL1H/Y�I���{�`txزrM���_7�:=Ri��j�Hd�QU��~���T]�p�ONNcbb��q�����b�֗M!P�H:�bS?
QTHr�G��q��#lKvZs�|���a}�9֚eE�$�9-����xJ����NE��h�[��Ye���Y ������-<��#�NX�-@\<H7|�\A FLaf|�k��ո�0��
d?������8tx�g��#"ʲ�c��A-���u R�l��67��j�:���~��};,n�a��o��UR�a6��0�(Ec�:��n�8t���%+�*�������GF��H�T�����fD)'1<<������wܨ\ߍ��$,Оf=c6�ڸR�Qy���qk���/��pI�z���H��i-c��ѱa��3����=lЀd���ѿ�#���12>a��6���C���~�޻���3�9�yf�ΡG�2`}�0w�Csl
�����{y��t'�g�l[|�+kN}KѻHw�V��&��u�)2�Wd�u�P���(�Yݪ郇��!XCĲ�@x-�����ƮW^D᧾��B?S�»!舁����	��H�8i`�_�_؞[t�Ԛc��������LCk���	m^���~RF��z�^?et�U\��--y��>�OG3�egB�k\�0����?�)C)�n�פ�� �@v�A���2�g��+��?���n֞��7����obK,���e-zoUb]/*�Dc���5��禙t��{��G��)N=�Z�ݤ9�V�n�L��0��(�e����a��*�J�=��U��B��t�D�O��t��!6�3��z�	��(�k�N���k霊�д�=��J}�UYx�|�6�46��Z�γ�������ꡲ�*rqUuKU���bn���嬵ҋl,1���Fec��|�&qt�vU����g0�o��K4�&�#U��^��*:hT��v�cn5��}�6��`�T�b��2��5�F��~t"`^=+	�di'T�:�"�+Cطw��)�9�3h�A���U�9�T�4|G}��[�����E�k�pF3���������i4�J��$�Nz�k�t����>�X3�4��A���ab��s0�Z����c��9�'	o�r�a�^�je���{����f�>\�3�x�� �?կgȡ��L�&'�n6��^ʋ�y䆧ip��B��,���������Khw7a�bi�,���Jx��Y�N�b�).���͐6*�'r����H�"����׾J�Z�Fm�ʌk��2�z��a�l���Ma�����+f�Z4N�6f@P��06RC}s��Mtþ��D�hSʪx�󌬥�n��+;����޸˘<*נjV��8�����ٳϝz��~�w��ܻs��o�g~��@�@�N�?j�Evff�c�X]�g6Ðd-�=�j뵕�#u}듩��q�xI�ٳ._�#�I�vR�ga;F�C�n�3�_s@ j��lʪf{�fp�� �I�Q�a��CZ�����0��	��t� f}7؎C�qi�i���0�MN`�<� ����#�O`��7���N����g����h}h�|�-�ׅM4x/^�X�̴7��6��nds��**k3���Ů�ui�|�TO���9V��w�>/��M<��{n���jy��6��5���L�U����G4���{�����;�j>�'��O)����gPLV�(il��>�Iu&4�t�����YS � �t�mI�vUI8э�2+�4�'�׽F�ݮ�֫aM����tZ�]��.�ۚJ��6 �s)t�Ȓ��v��5̣駍���琍3Klm#4�i��~���������Ul��J�F�QP�,0^���i9��IIm}��P��kR�\��s��R5��Q5:Cc�s=r�sA�F8i�,���T�W�x}9�9����ĴV�0t}yh�>�&7��}����[����~�Q0u�>�\����MOэ��Ԃ�_^0��χ(�Q��w���іeym��N�H�$�qYΝ�[ʗ���qQ�*%5�a�Pبm��#}R�$g�����`m�2o�m[���869��_?贱�����Sh�6���{�1^f�ǜ^�x�3آ��{h�@㱲'�~��j�k6����=�ͶQ��Vu�EO`C&�`;��V�?���uHx����?�/���(��e����� 6�-;Wļ���_	�ɨ�M?(��$�JW�t����l��w��	�R<\/-�t2���(FG'�P��X\�:tǎ7@K������U3좈,���Y����x��h��U�����21�U:�7�e�QƫQ+!��^_�Mc��A3��`M���V�]Q����L���S/�O��O�ޏ~d��ϝ:mk�6��t֙�=����������p�7c#o2��0�F�}:�֤A��KZ��F��3�k��v����J��n��I>�� * ����m,y֟v�a��{�RF�4pc@g��֤��P�n[�:ǌ���.�k{���'�~�=���������
-cj1��I����Ø8q�X���>�^�/���{g�p�"3�$�^;��_�?�רY�?����B�����&|f�CG���-���)�������l9-pR�Y{�M�\�7�N���#��7p�Ko ?6�0�ǽO.`�{C7^o��Y�%VAn�Y_q�=���'�w��(��(..��h{G����B��7=����,PP��G�r���1:fo#�N��s��Fifv�`��5��. ����l;ã�s�c��}���h�����[h�=A������O�"q�0�^;[<#wo��Ga���+Ѵ@.{�E4�� �\��ƥ�&��w}$=�����yd��\"0ѿ��#<ρV�]��م�{
@%1���m��N�	��m:KQ#��$�n�ڵ�`���G��u<*n8z�D<m4��s汨EV�����0���g�(��cX�щ	ܽ{�X�]$� �����!��q�,}ܺ}�8����SA͗.?7#`^����f�,X�s�Ū�/E=-�+��v-"�bPU���U[K�{r�޽(3��U��i���5`^�_��3-U�$m�r�A�6�&�BaRF��:�U"�c���	{MSN�!*9X�o�vt{c��18jr���p�ٞ�b���R�������
��r�^�;�wc�j�M�f*%�q-�9�!�������^����������B�iФ�&7'2 Lq3�� g8x~�R%LѨ*(�"�mrE�c<��D ��#:�0�k�tjj
���l�`�Q}}g�J�b�K� �L섆'sc1���1��)XQ+A�o��`iO�pE�]fA�LʮY ɥ���,?`xSFb�|��ݻq��FǢf�_�3��ǬD�ϱ��G��n�f��Y��,���jE�,D�#�ͺk�j���r޶�U#�~ԃ e��wG�P�2�Bo��0�q����h�Q|Hg��P��#��W�l��9�}:Ӱ�5�;�6VN"������_����.�Ì!{�0��X�0�����͢�c8p-j�$d�����|�]�Gvc�k_A��_F
()��Q�\�����
��$�Y,bE�W�Ac����2N��_Alr�mD����ha���@��a～,��3��'��iz�'��,��$�$����ֺ��W���j����u�^�]%kk�Z.�Ub�D0� H�0 �&O�t�'����������k�)��=�'|��{��>OOr�jPhm��]nI{yO�X�< ��O�N�pkE��󲳲%� ��O��矕�s��1�k����o�������.�Jx��~�w�:6"���5���w��_���xW�����������7R`ż���b�����R�{R��|��{�:3���Zϊw����f́|��<�Ͽ.��I=H���,mʊ�&��<2a�ld���z�&U�Gj�{/vS-(����g?;^E+�F�{����F�`Vqc]�k���n�W�!�#�f)���G�Bu�j�T����i�����9�2�.q7�r�o8�0�/T��@1�=�UC��ݍM��yJ�xk6�
d~A%D&�{��E�1u�|������>P�D ��́�<6���Ԩ0�	L�`�����s�)��6�P@2E�˒�x�ۈ�Q�)[1�$w.��ϋ���05���6@ ��;�]�s6)Х�T9~�6�?f迢���C�%QV�D(�6���랚�Q�e�6�]hk��\��}o8&���Q&�E�	f+"Y���3#�A���#�V��t�BP�V�8'N �}!F�~0t�t�n�{0�1*�1�D_Y3Zd��8ǆfi�	iT	T I}�^fdk�5�E�}@5�c����5���y�q����c? �Z�=��"��.AK���}Ov���͑ԂJ�t[�[R�nXH����X�L�-c�J��Df$�Hq�����m��| J�9�FFu9fn�=����3�ͻ>�t����4��\�`��:�)Ikꀃ��Bd���qi����kU�x{u�#M�ݖ4nޑ�k[���O���sO�@��\�j0s2�-���5��=
R�����ڲ��ٓ����46�GHAcٓJٗ�ӏH��rI��f�BE&5�^�sG����$g4��~�A9s����ǲ35/7����PM�|��%������I��N����`��\[�iO#�bMR(�i��jJIϥ�G�f�W߾&剃R}�S�OJK�Q�&u43���;��՗�< ��%	8"qmDvomJN���ܸ�?����4WVd�6!I��z�����m}�Lp��9)�3��a'�Hr����/����<�舩5������ള��!�A�F-3��ps�PX�w)�~Xv�,��4Ϊ]����;��/z�?�\�ʢ:x���<��ě��tX`�q[i {Zfn�N���b��ATB*�n�*Fh̖]�Q�� ���?{��(B�W�Lt��w	���T�L�������ka[���6�rV�|��M�!M-�r���崂#���c�j��7�V �yn��8(켈��}\aZt�w���
�/��ǡ��q�7�Ӵ��ƌ���DU�S��ȞԱ�3�wr�K�#肣\ĕ�đ2��콄�1�Ơ������A���nXPj�Ò�s�h^.O#�M�F�8��6���G���0o�'w��{��!p
	���Z]ά��=n#��}��`-*CY 3#щeg{�
JE 9�m^�L����Nk\���wn3R�%���	*�2��3��$!	���C=uj�%7(o��o@� ��{����U�'{$�@��>bV���w�u�VG�����uv^{K�?��:��ґ;���>Y|�c�}�)���+z=�h�KO��:Z�q�̳��+�ya|M�T�����[A�/r
���| �~@��s�UCx��W���k2_����R��+G5�+�`��Xww{OB͸���O�ؑ��+V玪P?jS�ƫ�u)%��L��^k[�R]3�@�.�&��'S����tY�8,���g��s?~U�n$�3k2�����sR"*A��)��y�n�����Ͼ!����|��_����>|Br�f��k���7T'U/LB&Dڍ��U�� �+�%���T��҅���������a�Ŀ���fg��F~�g.qYmU�hY�����e���rsM47��:&\�,h������j�m���än��:��*9&���,�j��G'� >f@����W$GA%��C���֠k)Qƕ@L�n�@��"���ZB�wh��҉�q?�	��&�#&y\��.��M̥���F�dDN)��c�Q�ηtm�;��;���d�,�[u����h��gcU�\n��G�\1��q\�(�����euu]���/����.a=1>==+��;NC��B�a����Ӧ�\�;�&����S`<��y�d�a,J�k�%D6�X�®,ևF�A�R�$w����C�ò� N�2�*i/卶��6�w�`(�ƶ��w7"P8�g��X��:�E�1���*-�Ũ��S�`�̏��n��f�$�X��2���r�#����ܰhl�ZR?^���8�R�mZ�3%�U�gd�(�Qї��5Ƣ����
U4HH�a��I�bseJo��i�W�T������d��v��O�j���i���<f���96�:�_m�N|!W*p� ��l��#B���݌!:�pΕ�PB��g!r�_Rr�V��zC^�3r
�u��Omn\�����'�?{M>��ϫ���&����'���嶞�NG�ӓ^�(�}R|h��������XAZ�=��d����^Rc~�Gg8!����7~&��Qu�4VK4XТ�sE����Z�r�er����~Αy�u�
�U1r嫡�XbgyU��w)��~�U9��-�`K�oI�ؗh� �������vD^y�y��<7�k�x��6��Jcy����,е;^�͞����ܔ��]) c���؜D}�[Z�믿!�>���A���99��%�������H����>��,�#�eÆ�p�ǁ�v��S�?�y���ԧ�EW!���jP�_�En�j$8hԈc��ys���<��-C7r��}� &�T�z�L}=�Q��#3��٧�����ovꌬ���DiC�)�^\�6n���܇��(�3���!e����tavej*�24����s�f�a����BIf5k�a\2@��8��V��<���ղ�����=�<���9�{'QU�nvNU�nݔ��ۜG	A����@	-P+ع
��z�h�!�l-Ҕ��#�. c���a���ӖKhrfd:��F[�!p�?���$�L-P�O�����]IM��$�u����{��w�I���Č�: ��u� T������S�l�2�cB�E���; ȫ�(�~S�n���1�剕���[(��(�
E+]E�M�D�3�.��'�ґqg3��Hc�lc!(�<�dнB�l�m���(znyg��&V"����S�n�DP��f�U7tmdT#�	��ޖv��haP�9i�c0p�@���А����a���������x`��Il#.�OW�lDi��Y�g�O!I���$)�d�b8����	?�vj��kr��u)����2��:*iJZ�I�LX�1�c9yPƏ�g���C�-��"���C���hzLv�n@��� @3�F�պl_�,#O<*�����/~N��'%��H�����Gߒ�xWj�~���|�&��Yi���ҋrF��Ohy���h@�N^�]�)��������2^�nX��/2s�����g���e98��XK
�)�16�\��~S��˗�W�Ho�#'�KK�^�MC��&�C:��l��q	�����ӱ#zmN��$��ْ\Z���Q)�=�����ܼyN&�>%G:!_���fpR�ts[gߔ�溾��A������2�����H��/�r�'���]�3��d}�,�v�ڕɑ���^�lv��X�F����d�˚=�5�kw�������
��t�0�N]' �DpS��FՍ��e�BM��e_�3�<H��юk�N���)mEf������C�nBR �9)< o�G�CM� [��O�A\ ^�8�U!=�;����H�R@%e�v�����<��b4ȸ�*���`���[ G�c ��70������x��{m�L�6 ? 󛃘�Y�O��I�/��q�h0i�!{	��|�/��ơ�l�wF�UP�"Aɝ�1p�i�9T�[��4����pj����cl7�\I���Y4L�n��u��v%����ec�����n08-F����"�w�k�j1c�3�Q����ivZM���!�ȪB��]�ߘ1�A���d.� �G��s�|^V���6���p�{͆��/R���E���׳�I��p8|O�z�0&��an�T�kY��~�� ʓ $+��xNh ���1�W} ft�jhA��i�J��Z�����==R;I���S�Đ��_�-�c򗧍����߽%��7dL�{e���y�)�IsS��HF�T�vd���2���Oڬ֠#���~Wg��y��?�1��YM��4J�͖T���}��N�'u���9]3�u��LU�z"+w���|U��Ψ�+ɼ:�Sj�7WWd��?����R]\��>�kT���W�z��7/I��ɤ ���:c8�=���%=�������H�m�ڋ/���e�F��k2x��<!G��R82Ϲ�jtD����k��V�(x3�夼��T�'鮮�v$5��C�=.�����W�wve��8h�H��+�o����i)>�~�� �����|(Ә#���m��WϤx�����������a��u��,!��e�Zt� ����G���9�7wYi��{�^�"t�����U��Ԉ��D-�@U �KdǬ(�cA�.J��wL��oȖїF�^�t�M�1t� 2T^t�����'2y8����\&�g��5��;;�r�W��D��X�VtZ��#ks���Z�3+�[�����ikC8A�C�<�OUY��7V����g���SX3�����lAO���b���7�������Vu����&���a!�yz^9�BM&C�?��}���������$e4�����9��X����y�OS3��	y˴Q�2P�K1Nf���Q�9SL%g��p>(�x�b4Cw���=8��!rӷl���{9C0��˂g��q�HU���Y3�� ��I��|�!wcf�A��H�Q9ԫB�|����Г�F��qC!lV S�S�Y͘Q�D��ς�e<�*H��zD�ǎl`�X72(k�bF��
X5����e�����)�!�{�ic����Cm�_����B\�'��Z*���&��5I���!��N4�mK��~�$poܐ�ﾠ�S����8�;˲�gߖڍ��lh���\����Y�d���K��$�=!���������LhT.�e�%�|E?���u�����6��kl�;�g��ݒ1ʹ�w�Ɂn_UG$:{N��"�LMK�R���T@��R����d^�G���fS/�L��:�O=/�t]��5ٹpA��c���)��{�CY�뿒����k��IU�]^���%)7�$������D�ȫ�~(`<���D��t�\�ѻ��zr���H�y\�'�jzڗ����~"��+��κ��e���wdbM�?6�ʹtn�˝�$ch.�c������5���A��g�Lh��;@�/zdy깸�=5XrS,��^\�հ6nJ�f�3�Ub*j Tb�<5���(�\C�i��0x.{D@���
���й���N��!�k�X��S���9Y��MO��������|��/�#�8�AJy`H���ZD��ω���g��2�e�fvt���}�;�ℬ��s�s�$B�|����>a�䣶��ԡ|�gj?�~��Z����9�^b�ݏ�5ǎ�=a�����g�y!�d�:�4�l���0����de[���τ6y� ^��9��w��P���a1ψ� �J��~��d�(�SA�����=˚�A�C��k��\�CC�kR��D��zaX�g:2�ܠ+�~!8-����a���K�e?��9D�8��[}�Z���Q�f��)��n�oR��]z����!���M�iP�쀰�Ч9����5��n%w_�R��R0"`�B�3�� ߳����YF
��͢��F��~5?�*�W�HY��dj#n��6A{`��޹#��^��
2�9(�a���s�*�Uԋx��vV�b9UQGx[�㝫�����/U����5�6�eD,(mvZ���|�L j�$�qKJ$�ii�q�*}���Udvb���[/�Pno�"�d&5Cz`�.S�� Sf�������X��/I��hP��ѯm��@`�w9�&�����t�}W��A���p6eF��4�ݛ������m�S��������?��h�//�J�~����{^�J����Ҋ�4�� ����'�|�uYy� @忢��so�Ʋ�Ku�|E��jKn���>���� �P��	�~�(AŻg��#��X/+ǻ�mN]�{�Ğ�8V��p���N0 QŞ@��T���&��g��F�ss��c��߳@!��X6b�C��{<?������a��ay��G��� ��5�4�v#�ZY����}���OM9^�������؁�<h��6賯�s����W�]���&6�Ǩ4�]%զ�����#4�vM�a/?��y<Ε�����j���!�l�f9�G�?����Н�Ҩp��s	h#y�#�f�C\�vړ�[e�w���,w`J<�̡�%��p&Fb �		�;�q04��O��Ĕĵ�� "~����hW6�!�[���,gw��N=�6F�J��yz�!(*Q�B�d}���,ؕ��B���#�A?�&��H'KX��:P��x���b�`87+�d�1ʨ M:r�3v�9�l<*d}5>-�8�-��>�l�/I,@�嗏�Ġ"EO3vU"��8��:z_��JMOTiPRZ�s�+R�f4�A���;z�@�u,��,�:Q͊D���:�|/G �\_32]S�u{5��&�Pw�@)�/�3��M>��NK�qK3����2����=u�^�%��]����S��tQ���;5�!)�5.k&� e���nS��;R�PʪH]2����H�60j�D�A9��~FUp!A���J�E����Ђ�m� ��bݓ�BQ�7���������q����jƯA[;��W�@�S+i���ޑ]��=��,�W "���� �	��<�a���5��~���&Y���doz8�۔�m��!����Yz�:��0`��Zb�k�F�̩c=#���3lā�if�v���F\e��Y�L��V!���?I����Ϡ�ń��T�0��{@Us�Y$6��73r�s�>������5�]zW~�S�>�;���@�Ӕ������ ,L_�#yH:�W����[��$n�;����?q��7��8?0BX� �	���PG�K�w8���@\@s����ʡ�5�����\�.j��q�����`s ��ԅ��:r""�?FTMD���8�g,ދ3�Qo=2{v���"�E	������aoW7�#�9rn�%����ې�@��J�R�o�(�����z��W�F�����u� }�ѱ�FeW����,VV���I.u�����";'.�]l8":����}:,�р�6B�F訌�Z�C�h>��r@�ʇn�Vk�f�e?+ ��/ٕ8�. �^�1EGJh�EYЬW�:�Ts�t�� ���*����d�A�fr�����Ϙ}p=�N��mI�1�ʚ�j�	�i���%َ�$.���9�I��캭Y�>��mJ�2�@P�ѓ��kR&�aKzݖ����_�n1ӿ�s�z��p�Z���+�e�Gb?�X��rdT�NPL�u4��j��G�H�w�����`�]%D���F�4�����>srZ�sl�t66����L�����ﳃ�:h}���%�o]i���b�>_�X�O��ԁK�X�;=�1�'lb�V'0��� G6!�,s�Px���HO8v -8# ?���X�X=Ƅ�@����	�!��M�K��7(|nd6'=�|�� �N���C��(�
8���}�Jee��fϴ7� �''&ecu����@v-vٹe�Ƒ�����>x;`?�9~�����U���D�8�*Ć����[��3] ܈��Ӟ����;KR�V�������Sa�V�cv���aC�p,�X�b�O�쾄��#(ۈ,�]6��qB�!%Ż_���g:�n����=�В�+ɐ����.�r�����2>��\�����H:眨8�-eW1?��&g��>K�@kc�~�fNQ�.�ݑ�:W��J�C��=�>�}zbar�Ƴ>:Jd|�Ro{��q��i2�u���%���#�k������U"�����1�{"T#��qc�csat,�F̬�m^��OI� �s8�!K��f��&��G��8t���0e$�T��7��J��Op]�=���0f����|pq9<��  �������;'}�� ��|�i-�y^�"(B�GĄ-�R��_�Hs����bMxsh��+�H��KtrA��Oh���s�9�:�ɢ���y@r5_��(L�@^�P��ͷ%���hA�'55^�����i�@3_���b^�I(�RU&O����4�M��J�X[�/��߹RBq����d�7eD���Đ�w޷@K�)�	,.��C^ίs�����{sS�;�(��>+�<�#����*��ޕ���T��+2�i�\Pe��:2x�؃v}$e��1��b=��@/ N�	 '��d�y��=�E�i(� `�~{���{������w���mO|1򲇡���
�`[lB=Љ����{����i�{��Y�>cSD���4xΕ+���k�!�FF�ޜVL���pi�3���h��J�^#���6��S�WQ��p�mJ;+�����ȞMM-���/�{ǝ���>v�$`]:�����fӀS�2�?V�մv�k�F��B��*b�=c��2ط6`Ha���Z�{#�J|�z@�J��S����V�����o�mT.����f�Ń�f�9����+���s>����vX�B�_.�H�o|�@�s���>�6 [
����і�!��Ȅ���db�P���"��Ɨ�������
)mL�������c���z�K�	����$�9G��l|�F9���F�lF�z��V�`�76��k��&z�M�N�Ad����.1G�Rn�M!>��ҋa`�
�Y���ą��qx��"@��#��!��1d= �Ab����h�vc�BM��4��c,�0q\ޮ}�S�<�����-���s�C�`1������Kd�2����9�!�E�_cD0���=];]WM�(G��5	?�k�m��#�,S	P�N��]�t�S5Z�����_�|GRur��� f���>�eX�����*�L˩���T>���<�ʧ. r��V��rV*��O������f�%]�N�*-&-L���O��Zh�l�r�3>.3��%���sR<pP숞_�Y�ڢ�'OK��G�����~�mA�x��(��.s�QD�Z�'�=�9�(��\V�,�D ��0q�V��U��~�Ꜫ5ZR�z�����}C���X)3o��Yl�Z�0W���I�����禎a�>!�Ll���2��_�{j�z����MϧV��%u�s�8���@���_!��$�H[B&T���:��Z0���e�4��SF�i�G�(v�|�"[mFQ+�����J���� 	�<�i��~P�d|�X_�G�p-=7E��k�u������g��<�����µ�AzU_�V'�`S7�D��(  ��li|��(�M!�������J���L�/Ǖ����?f迊Δ�{�峦w��K�4i�yI�M	��0#�X�+�ʺ��,�~_�J�E;h8a�Kn�FF�`���ƧT��d�~�?5�1���h���9�FK�����4�X��Ek$\�lNjO��(Y)�2�Q�;;;K�c Ѱ!Ћ"*4�qA�N�c)Y�6i	��4�.c�<�EY1���.�dЛ��&G22<-��G�v���noʘ�7t�dc.���A��3�G�Z��,pS����S� �W��#��A��"�R�62�~K7�j�!b�:j����=��2B��Pi-�T�f)8�(�g=ל>PzG��!8��dL��x�
/�Gg�l%�����[�JO30�Z�5؃�:���y����H���j_Z�4�����@�l�� ��]Izh�n�8a_q�Ej@ӱ1��Iu��uMt� ��u0��f�a�R^�
��quZ�i<��W�F����/tΙ�%}��bf��R����?.S���ȩ���� �������������Ž���X� 1�"������z�\����Y�djx6k�9���yY[*4G��u�m���YP����²fk/��9ǯ$!y�m�������x�bA�ib��75|����;���: ��欶�N������7��4�+A�O��b�<s�����j������nnm20˻�;0�T}}Y{�͂�<�|ȳf�~�=]�!O�'"�S���C��Դ�@cR�6�{�~` �HK`�����#?|��� p��F�����j�hW8:D�~�Z]��<* 6"l��>�%����7�S}m�ߣ�Şlc�";0GY�\M���S���ޣ�&_5̳�b��Y��1C��|8�Ln���n�����F���kX�4�	o|}t���������7%x(��=p`���&�#*5���J�f0DINy:l g�c��-��9ޡF�wޖ��y�����;1>I4j��%��P��O����aJ�d1��#F�
�ǉ�=29��a~����Yt�=^���`u�w��yZ=p�*��mvT7����D�w�%cm�JmC O>�Fm|��$����P|���$'�#jow7�2;�Ư�����Ȳ	���і =��W��0:�� �3�0�(�F&��캱�9������q�	�0�χ�?��{F�-!��.f�#�̾g�
�����ٷ6:�F��E���뤦�L>�4��p[G�s^���>5����Z��>34�n̒9VȠ'��$�IH$fH}rT0"4�m��6B�
�I3(�M0����O|J��'�� �,zx1��+�����Oʑ�7dy�;�ǌ�& ��gmբ���XD���~�"������I�x�nqz��{�ʩ#zI-]��:�{�{���"���5��j7��Խ[���J�gb(`x�>B�k�3��.�'��&�.1�hh��<�004ak�6:�@
�^'�*jB�M�9�|�
�X�#(`[�����}%��:�28��;J�=�$ɉ�ܨ���b$�R�@jU���`=mT��J��,{vn� ]��= � ����J��DX��f���&m+��x�f�ZN�-
L�F�ž?Dx|�� �!8u���{�?9(2j��5� �wd@�����)=f8� '�����r�p�i�����°�����xݽ=��4bi칽n��ԋ����-5zAd��5v#"d�<���Y��5�)�%� N��l���!�N9M�������_��Z<*ss�2R[�Yf����� 	�@]��h�@��[��)S��+�e�Gi�zX�B�q��܆��hơ?C�������DԿ�F�����T�aV�9 ��aXv��u�4������60��9"`��F��� �X	N�C��64��5c�Sz��3�C��ʧ�ko�J�:��&��L?dEX�e�]��Lpߙ�����E�g੏�>��_��|� 9��RD(c�
�
��,��
��{x�XU��\ͣSڧ��^�ᘺ�\����%�u�q�dx�(�b���Ĝl��YrMԝ�ƺ�3���c�X!"�0�M�Бaj��ߏ;,����ִIϫ�Dۃ�:x���X��G�ݳo�އWI��)���d�n�rd�I`�-q���ȕ����]�{��a��^D�=��s�ٛ���r�&����=O�eG�3)���� j�w���ZCk%P��Xk�W��,l����.�x��ʕ8������c���@+n������s�m#���=7:6���T�=i8�i��;�~zbbR3�m�`~zĳ�C����h%}��Б�d{ܢi��A���4QA Q�k��R�2�s��+/��Ԕ|��P��$�<*AVAL4ؐ��5N�p�9���n�Ԓ%������1y�y�������L�Ć^猿�VJ���|��#����k	�C��8�����դlz�>x�7��`�cv� ��M4ӛ��59ʍ�~����')�B7�<��-a��� <��ɻq,| �n7�)��F� �r�f���~����;w(3�>r@���M}��q���E�q�,�]�ͱ'��S�1��������{m�z�*G�!�����ʀ���6����.
����+�L�͗:Qq��jXvu�D�OX0&7T�NNa�\Y�=7�v��rc��`d��1��6n����ãC��<�'D��g��\����O�%� ���@;��qͭ]��`�r�9y��<�|�����	z�z�ܞ}ݛ����~�/���G`_�v�~-����S3t�fn�/���22"���R�ZjvHCdp`�:��@����k�A� ����R(z7��6&�x���S>o����4����Gp�~��H�3Ǌ���(����;zD4ڒH�;���BΖ�ow%B�2X���,�:�H�v�!7t�C���B�@gFR�fp)�����殪�ٞ+�����G���?;wnAF�BOm�35A���!Ȍb��#�Q�˨q��$�
%j�Y�A��Z�P��E�>/䭺��]�,e�|�������VAhj�q��]9�;@��{n⾐P�"r*�(i#!�q�:g�kd�3>zܯr�F���t�	E� 8$�|0�_�])�8H�{${���,ؠ���o�����������z���	�HJ]�2�td�x=l��+�9�!�$Q�JP��TN>gjtH���F���ɫmi�lP�P����������fb������t���N��=��7���#P��q���COl�23�}��Y�jK��Z.��Hk�:c�N#0NX2���ѐ�����T(� �ūP���̇9�^}s���E�}�ȡ)�>J�y�|��;}Z&�����Q�LuV�����g_gI��[oX��3O�����I"Y�U���1�a�X���ܼ)�YEa�����v�$�� B�Aq,������m���mu�{z��,�C]��r=�
78N�{��ef̌A� ���=�H�0��)�q��|6]��~�Y$�w�H����bM�ʥ��K� �]͆
��HF�k�?u"9�V���a�=Gja��x�C�����?���c���A�
���:�*�D虣ثz���q��s���M����Ꭱ�7T��Z#K�(�����kՁ��Ը�F�i��Gt �����?�>��i�IY�|� �pں^S�]d��z�xPYȣ���R	�	Z�z�3�a�#�L�l!W:����$g"��EƖlok��<�x��R^I��g`2n�:k�������9����q���N3`\�&>85�kf�z���vS:�
Ւ�3}�����4��ϠE&��'m5��m;7�J0���fm.싾k��������7���ɬ&ސ��0���<�.����2�9�w�vYH�X���M�:�z����]Kϧ�A��I���n����
������W, ��y�,>2e9s��8��{�an2�Z�9M� D��U+ �V��DcЮ���^������Z��a �\E�������v0��jBso[|TC��4X�K�\:��V��w5��b���~���C�1������@n��S��A>Q��� r�Dΐ#D��~T1g�,*5��|H�G���hK�e���:�,2�B������]-k4���)��S�W�±P(�g���=zL>8�>Q�ϩ#��w��s�䓟��<������.9u9]��-�n�t7���Yƽ����Q�L�2��c#���g���!(8�� �Q��������
���(����1��2�F�^Vc�����(%y�hx��|`�jv�cFYePև�B���0l��,�k�oq$��Y9���8���<�t�(�Ѵ�'Q��D5�C�/��ڽv��{Cc�=�{����z�~^���7�sT�W�t~�6�zÉ9t�6�Ş���x�������B=���h���sD�rV�����}h��AL
�X���H��۸��J��;I��V�#�f� (J�g���Ñ' ����ɪ�~^�B�@�'a��:��� �
�'���CʩV��&�V%�-˼S�@Y]��d��� �jCVu��dN�%�~������M\��G�|Yn�e�N �v �[�+η�6�p|�0	�O!8��U�w��@+z����iB�9���7�P[+��Y�A!��y�X]�ɹ��N}wsK&�f�9z%[�*��hYcuT�o��$���_wW�$zוZEmV����ĘrN>�U�H���}j�Qi<`�\��s���N��Y�X_�5���m�w�6��
N_Dr@��{{����`h��:ݻw��u*ԡ
[I�{E�|��U���j����=ϵ��b�
��ou����� hjz��
���-��e=��=i�mJW������A��N<?��I��r_<���?���K���Wzsr�����^�����I��fs��]	��d�1%q�Ն�؅ԁ�Z���dq��g/��j� ��܌/�78��.H̜Pse�lmnȔf�/�wAf�r������:�B޸y��'���8��Ϟ�o��_h���<��C��vA�HG�9�:�`C�����c��D?;q��8N�j�VW�i��<99)�z�hս�6�hi�|�v���#/��G��k�B�`>g�h��Y_]�ջweM���^�Hxx9�G�l�lw09z(}ʾr }���� b�M__R��~�n�((j�+2��VB�5�ݵ5���1�IA�"Fy|C""覑d#�D���4��[	9fi�B=�]n� �̯2@�d w��k ���2H��ա�����=N4�+8�%��= �`\�7�1����5���aN=�^��Z�H9,�Ich�-� �Ɛ��cN�V���I��u�]�Cv5�^��E����@.�X�o�וB���
�㡴ћ��Om��m��NO6��^�.���[��7ޗ�r]O����)v�"�t\��-�����i���[�>�o�e�u�u(9����@��9�#��BU���Ԯ9����+LM	щ��PIP\�@�:6@p�d(^1��:a ��x�oޒ�ӧeG���C�!�7e�i9xpAĺ:��˃���Us��¹�//y������M�@^��18���<������GdY�酷ߕ��&�U�?rp�p�ǎ�s��c_�v�f�s�eK3�w�]�d3^Q�5Ͱ�v�9��RxKE=:��m��u���.m�^�� ���c���*ׯ_��X'{&&[r_��?�]]���G�/_��sm���#�����7��6�z�3�>��Z�BZ���D!�l��5���w@j%b��)�#�!�6�R����:��6c��jQ��w��u�Ӽ�z��pKW�Z�kh��Ap��?��}���`��@MD�������t��N����9+!5H��� okV�x��0��6��I�D���=GҒ�A �B԰m�_�zENܺ%'�<�����h��"XЇ�O�����Ki����?.�N������rwyY#�z���K9�����qѣ�m%�p���j�Ǆ�UO��Ѥ�ߕͭ5Θl�6f�2o����ɓg���{s{WN�q�ܞILnk���O_QC�,��1�\Fm�Ϸ�e�,��P�1J��{���z��� ��Fl��2{���$�{�Fc}m�e�vcWjPB�>�����熾g��z��-���|���	�=ǟ}o����N�yׯE����~��_�G�>T����wԨ�"�td��`�9`�@{�@"��Q	��_����V���~Rs Wb/���э�2�(�=h�4@�{��u��OߐW��]�7�e\3��f?��xT���rx�3�hEA�πbj(�xc�/a�ec:�J�}颌?�Nە51����ge��U9�� _��W���CRVc�zQ2��tH��9@TX�GU	m �[��}̥y���v�C��)�Ơ�sΞ%�{�����02s��u��EE�M�:z͎��ҽ��1�=$ �~�ҕ�:���Bl~�jA�>j���,�w�k�E�&���أ �5:;r��r��)9��[�Ȇ11�19Z{���갮|x��w�5b�u�:�Oa#vvw�wv������-v�}����� �ժU�.-ݾ%�����|D�K�ɷ"�s玔4�������6U��p�ֳ�
��^xA��봙�7 ��lG�ۂ�R�ܨ��}F�Z�ĂXW�C��i �{8w`�,�.	�_�~m@,�ՕH��j6�Z��m&9c���W��^j�Fqz�MI��^�w*VC�׈:��<լ-���_��i���������>����0��P#Sp�ݸ�m8#N�c2}�p�]~___��7o��d�(�؁��
B��Ҍ���~��<��#�}M�<����|�D-+���G�9�6�M��Y�2R�L�Y�y�s�{�`,E?�BG�������y?v��U��W�5��Sl|-V����rQ����RB �! �3��}<(��^9��n8u�$l�H�<*�`�G�TJ tAy�< �>�0�M��XU��]��9�;���5���}t�}�UM��7Հʀ眚�o߹��D�e��.�cw�ApP��-5~}8��*b�����{��ݐ�f?# s�
R��f1'_����G���q67w��!,�?5@��O��w�S:��$_��C�����ɛ�=�k����~]J ._�*7.^��Σ���R����:t�/�4��1�An�9�^A��A1b��ϩSే8�q��y�ߑo���CN�<.�~��2w���Fǘ��DǺ>w�`��)����`��A���X�o�>)����b�T�K� 9��.oCJt:A|����^J"����e�OSg]d{�����%	�\묱�-��1����h���֖�Y���G*,u'qA�b��.���
A��a�G��x��龫�F�"���2������7d�[[�2R��&0^��_�DP�%��l�l��f� *R�8]�-�j�n-�l_ P��ݾ}�	z�-d���4�������ޓyM�&�g�$��K������9�h�<?�>�d����٨��b�9�̦�����T�8���4|��G�Z�kn�x}$9]�U��^ׄ.F��ܲ��.'9������~x�W�N%�<�*[;�(���v���R��\�͗NOs$'��MLM�Ｕ���:bC��@I!�ޑm�Ĵё9Y/5�JȦ��AT�)��VG&�T(�b_f�zТO����(F�67׉-g���X?!_�җ��˺)����d��U9�����rT2�V���纴�$+�A!�h6��r�G��\X׍�K�iʮF�O�<)ǎ���m�&O�>�*7�n��۷ա��Q���"�,%�T�;e4��"����ٿK���'���� ��m�Xb�=x�LWH;n޸&k+w4��,coS�VC�(��W�gVF�������P�b�HxTF�! ���9cI��w�f$2���B~4C�UK?t���ɺ(������ʷ�+#͖����b�E��ή"wK���Z���c�K}l��u�Ea2 �PJb��b��^�5T�V�ؑ/]�,ݝ]���{2vl^�aL�������\�+��q�_�$SМ�e���/j�Y�����,�>t�B�a�06�P��Dz���r�r�Ă��@����'���kr��O�3���d��)��Qb��}P(�O�]�ީ� ϡ��}�+I7,�ZK�T}M���f�]�έ��;����2Jn8O�u�VQ�n��K=G.�(-��B��kT����޺%�3�1vȈ�fcq�,����(K�,����ut2�`'g�Y�9d��A�D6��@����yp�il�kY|��9��dd&�� nh�a@��C��h��=9>6"��cD��Z�� tT� �꺇#C��e�X�9������p� /qǆ��o ���ԴM�,�Y�k����� �F7�_�"?y�%�4�F�;8�g:�ḍ���oh��g���쎏�{��g{�M��d]��و����� /��d@���nSF+uO�v�y�ۉ��^�R�X��������q_9����7���Ş�F]���p��U�4C�C�'0 H@�x,��Q9v�lj$��1���-�
IP�^��\(�Y�A� �@���o��[����]J	�L�������;�2z����A�O�F� ��#�����%��������L�L�u�$������M9rd^>��>VP꼨�����yO#cl��h�����G��$l8�f�JQ��c汾��@�����q:s�����;uF�f���&�Y~��w��w��o �U�>+����_�d�CG|ùV��s��G��#r��lʋ3�����f������H��s�\�+0})�ԇ�_�89cD�an����'��0E=C��v���}��&�w3�F�Q=.���?҇G����m� � �y�ӟ��N��*���ve�G?���/���=%c�Au5����u��3�Z� ?�*o��@F�#i������mM�OPPg����8��ܸ���Ԝu%�L.�!S��s'0*�<�N�I���j5Ѳ����@!�����|�?���xD/,ʔ�w���'������;��OM @�. 
�r���X��k�ѽ���hY~��A�����7�����}GR�(%��seY�#j�;�[Vk!Qݎ��7����
a:��Z��P�ˎ:ߛ���'t�ݹ#������(�Q3��5����b�m�f���,�~;�XJ.�,h���b����{�qm��hgvw��R��]�ܗ_|Q>��ߐ��I.Fx3zOoc�Um��C���,����;zX��(G`3�[̆5H�]����)Z9(Y�t��P`�z��&(������*�� ������{�9�+��?��OV��z�$y^m��H��~@P�
 �a ����92L�B��'6��e��ө���b��	����9��|dҮ�H �����%��w69�|�c�����5 Y��� B�O��x�W.fЇz>�j�������=��kI7�ģ�ІD,+�T-�:գ?"7nݐ��و�I��9�� ���KC�6����6ҍ�G��Q%�<�k���(��.��؜\�vUr/��矑��4FMۚU#
���?/����n�0�MMɖn�-u�_�����C�u}�ٙY���a�p���!�;�LHl�c��R`�^f������\7�WՉ���z�O<�$��FcMf��ԴqX��{G_����Q��N$&�o����m�1&5��,\�2JL���yP,�SG2�xD..�]�/ݾ!���4�z`nRڕ����;RC	T߻'Q�<�~*Ó�ת4 �ӣ��9�ؕ�aH���D}o�b�e
YP���3�+s��Zs�*d�Cf�p���I����y��nH�PE|�YY��g$X�3'�&��Yv����5����cy��'�������Z"w6e�5�Ƈ��\�y��e��-�6��z�b \ÕA "4PnC<���'���a\g�gx��7V�J��������D��J鎬~����dZ���S�O~勒C�=�p*�Jxq!�T���vo�������Y��y�8-��w�R
'�ʑ�ޔ���e���Sd�0�,G��Rln_>��?�K#������kbV��>�R��nb�_(�^� ���hG����2�4ʳ����o�X��u;V�����Ae#y)߿�N}����QUp`Y/�4ph�:�R�8���x��|�YY��&&�)���jޙ�$F���~&�cl�4Z���0�a�7 H-d��F��KOG��DJ�2u�AX�Y 9�#���f�Ǐ*n�s��ɶڒ��~Z9�7h��ߟ={�|H�H����V�Ȉ^����t\	��b���\!�EN�XR�b�������)��{�ɏ;E:��A��X�u[v�7�6 �NZ.�Wu�/{�|�����g��}�Э�����-���K?:��l����tA�1	�ဢ3�@&&'�w�k�Ա7��@	�E���PӖnt,�CЁ�n�ZQ�'5"���o��D4�Ʈ6��w4�m˗��%�W��J��W5�����_��LL���~�r��FD��O�\�z�IyX�:�27;�L�Ν%7�\�9e�|�e�4��&�jև�ͭ���X�iZ���?����a��eB�����C&�_������+�\/k��I��
^�3��л�⁕�d�h�xr��(�섰8,���A ҋ����FG�������|]���^�ёI9}��\�iɪa#�dJQ"%�j�3X��ԯ��9Es�hŀ��h0b�^�_��r��G�H �IM(7�x��G.2�{THEW�u��/�����~A���l$j`��rD�՝���΅�������⿑���x�,��O)STmF��!`��ThB�X���J1J�^c��1�����6�؊|�Oě��N��ٕ)��zN�1�!��E=�k��PՑ �QC�w������f�{�z��\ۖ���޽%{wnKe�(������O<�����lh���8�>a��ʎ��Ml����u��q�����R|�cz����g�9]sg���%�jJ^Sݲ����1�u����&�/Ab�vjc��ЉI��qG�P����������ۯ�&�����D�	��\I�;�o��ʡ����+��"L�aY'�{=ض���,#X� ��6���" �{}��$���>��0�����hP���u)$�Oɭ�y�q�C~&��+X� ���ځHf�v�ނ8���s�I���YUD�$�#A^&  ��IDATgÁ_(�h78���\�Eb��G�j�|H�p]�:/]����U=a�ѓ����r��kdD�/�Ba6�6��c-3#@��=ɩ�Q;���@�{�*���3���Z^�H����]�M�*\���G�+o5��.�� (�b��c��+�Pg��Z#�؋6� ����Z�=u�	��dE���L�F�P�^ZY��Y�m�pdo�N�#f�`�A#�6�T��^��f��4��ݕu�<2ru�����qu���\�����<�Y�ʰ�j��r��M�m��g��G�xR^~�ey��?&Zu��y�G���w�3���m=�'R��|��,����Sy��TK6W�ا�}K
��j�$'O����)1������!���k���}^ΩQkk�Y�T|]� o�^@%'���Ei\Q��dH���dl���_GFՍ[D�a^6-ξ?��s��/�uN���\��T��X��d{K������1��4I��DB��jb63��Pߵ���@�	#��r]��3�����@3��f]��'`����Г�����H�2?,H�3�T�{��.����8W����k��s�-^�O��?����RǨ]K���?�$2>:"m̀�(��j?�7/Ǻ���T����`��,�?����Qǭ�O^~���-�S-�F�2�Y�����qcA$�X���Z�+J��8���e=WO�U�k��������$;;r��y���3;}XB��A�cd*�a�/ tS��{Af?�h�6X��5�?�(���{2���d��5��tM���2��s�߹?��R�c)c��)nA�� '��\��m�9p�t`�O$����z� 8dKk�?T��z�oʵ��D�/_";ޘ�ࡨOV��{�	�?�(7n\VZ���њf{(e#6&	ڀ:��f�t�ibz�D�<��Y+*�w��E��҅�LN�~P���]���cd��� ���NPܸvE����"�<��H��hi�f�ŵ<8��QҤ�캃�6��;l*�ח+ESg>9=�j�@�������G�dh����+�����+�Jt{2е�*�$X5�C�=�h�'�c���&�)���� q��`;��	���Q[�t=�����@U�䱣R�hF)�ʭk7�cO>(��e�n/qd-��#M��n*g�4�E�	#a�@���q�9t�3 ��H2
m�"��Ѡ1����ޑ��J��$���<|�H�;21!����> 
ܸ���JG3v"��rDV����0���g?�%!G���O"��k%���w�>��A����1��1rwu- @�ݽ��������o~󛲾�.��իWY*�'���X�z�"Q�yW�'�1��N��V�(���\nzlJ?����hJd[ꬫ�1�?tXf�N[[]�/]��?yIV5*�aoh��#&
���RG�a��ر��w��i,S�<��N��z򲶵%�=�q�;�@l��|��R:zP^{�%y��!y��)�Z��@yBI�,w�c{�ꄌ���L9?8�x!}��eͪ[���[���z[�v���4K�:� ��<���Ƌ�ȍ��!����:yɏ�ל�������lS�oO��j�%+�c�I��{�o�������b��E�����{We7�?Q�O}�dz��ɇ:�PR��C|���
�zV4И�W����'_��,v���2�����G����ޣ�5�ca�	��f�?�������gI�y��7����V7�`Yá�/�)]3?}BƎ�HqqB�<� Ru�R0�X�XE�Ѡ��ٕ��? �*�B+��i�m`t_>�կ��3z�Uٺ1���������g>!}Lڧ���_�c�C�X�X�u�(gh ��5�	��6y����5��8.����)	������e��-�^�&{��Ey�񧥵�-uT(�:����>&��y�(��/cݑ4%$�U\���o��&i_jm��4�7��aƬ��j�i����{���&{ۻ��S�ȸf���>��� �]�(-�#�͑!m��Y_[�;KwР2B�enE�ډ6ߞ���|�Ğ2}u`��T�8�vfjf��@�0#=��<��C����ͳg�ڠ��ui�C_]Y&�k��9M`w@���6�~|nC�"Ƅ�hG�4&�* �Gⰴ�,AU�����&Zr���[���z��7	��$a��%i���5o�I���z'��A>� 5�O������z`�M8��A?=/A�J7L'�A�ߺtY�/J�4'��,��"��� ���h�>ƅ�1��:<�N�gR�&�=Bi
�&�C���I���4�-����������ڈԉ��s}���"�x�qYX\��9�A���{�5���|�sT@��
�������|�󟗇Μ�s��g�?^
D�v�'�ʨ&���/�a���R�T##Y�RcEwW#�����@<BE'0N�{��\�����T�fa�F�a�'�:�km��H\l���R��q�"R�Z�D�9ʒ9���[�nl�5_��W������������/��f+��{W>r��O�A�\䞁��N&z�[tJ(!��L�N}B�e~�S�����zY��]MD�T���ߖ��R��P?ݑҩ#R?sR���.���x92~��<׫t\}}�&�;�a}�*��-̪�n�Nν����:�> �^]��,�g�]V����R�EEA��JD�38���������ΎHn�"���ý
��;EeluVF���#J~j&Y-i�1����\v�ו���X�U(� �E0�)��(J���nٚ�f���v{fM���ff�j�mOO�=�%�mY�$K�DJL"0g"�*Ǘ�s���+�Zv� �i�@�޻���w�>{����4�t	d"D@>��K���N�����[5X3qjI9'!e�#���,HzA��nNq�yL��:�<�R2b�����έX Q��W���?�����S��*�o鍊1��K�cHǚȢYY�,҂�>��:�E@����̠��j�7��F�ڤM���Xd���d�H�,�*"�&A[�oݍ��}B�ˢ�][��#AF�Z$m�4�:t���_S�����l�� �p0�ž2��(�ifjo���f�;n�-�j�2֭߼Y�W���$��;����9�9e����V�.+0cr*j��E�a��~0�µ��+�Fc�ŉ(���=/�O�iWw76H@A�yIq&���#(�� ������,��tw���v���RT��E�4Q,�mX��� -���(U-A�[�s� У}a�iI���Ś��$�����:v�}��9̜:���8=Zp[��t���e'�\�Eȯa�z�p������_�o��<�VX�s>�[pj[:��t��),ٺ��.eEjȦ։���˱q�&�#Ɩ���`vnZ�7�PL��f�ʗ��Q�#W�n�����"@H�4A5�TB"AӅf�(~ ���
a����8�޻�����v�Z��s�/�+R�P�,Q�����I}Hp
Q��s&Q�۷m��k@$�D�R;�#����"�;�}S�	R��ϨxL�����+ר"������(�	���z���&�|^gk9���c��g�2b��-�il�l�"80*j�\BfF�7"�R�#��5IC��\)��,~���7߉��^���O�,T�S�Q�����p4ex�v����]�^T�3J[r�@��s���D���T�ۼ[�7�^����6o��|W�뗡����2������Ā�ԡ�M\#�C�#�G������]��+�b�C;��JBS�"�����8 {���|)�v`����2�?�"��萸�C�:��2^�Ώ�p��vf����	�d�'d���+vo���0���"V�#փ�撱&ȍ@A� w4{Rdv,��֌dI������^� �������&R�~	�;֡��PU����Y+ 5��B��6?�2�w�,酧�V	�}�ؽa;���o�����ʅ��gy}�2L͌#U����@��t*�8j�|_&��H,ٺe���*C@0�!!�5O���zY�᜜�ӧ�I�X�0'=����aܴg7^>������D�&22�d+�^�1���]*��w(Bb�u� 1������V�P)	z�zǎDQ2�7�,A�tt��Dm�ٳ�%8�",�0*�uŪ�薬xffZy%Z*�b�d��9��q��'f�g�/G���kc���a�*�����*Ν>�N��<)r��=]���qUm:���産��q'��A"���̞w�'����6���B:-�F���DW��J�_�C�+0%k��ѝK`YW���AI��Uq$��zv<tٍگ8��@�K��@�v��:_��m�j���X�~��z�;��Ι���� .�R�'�R�(uQ��L�[�o��cGQ��`�6*�3��E���m�8E*�<B�
1,�FHYϒJ��C�ʡ*h?�(�*�^R�]�<E#���ב�q�s4� F�<8�ZU��S����>��-Jf1���J�n�z����#k�V���M[�	��h "�jt������ٍ��V")�}��:�%8��|�ǝ�ѻ�la7��d�,���`yX�L��2g�������p�`��ݞf��1Df���GT�c���z�*^޷_��>z�h�+9}Lt�S9u�̍N(:�d��Lc��rۇL���9�Ʃ�$-q���*r��i�Q�ĸ$����_E�8y���_�r���!��o7>��ǰ��_���Sh����`���iIA�[���)&Ė@(���F���o�/�*�&j��3h�К+!;ح)>K�FA�����R�y{1v�AMF�4�Y-�ۍ�1�T�kzW�W	�D?�tٓ�μfE���(,��J�0�3�,a� �cYY�ZU�r��g�435���{�"�QBID��#ڲ0-����;��=[̳̄��\�2[���Ѹ�ˏ��
n�u'��V�Cw~ox	���	�X\�E���Wށ�ƽ��Uݼ��=�3?}y�0�Qi�p�Qd���i���tI�⽀TI':\����O�S�4��\�D#gNbp�
�%�Kt�aIvG��Λv���wP&�&��
 �KM�칆���;eg�ِjyG�����4V�-�����!�i�K�杹NT%P<u�Έ�^��$�X�f������"/�;5rEq�!ӿQ=������9R��m�����I�T7�:#�^ՠ��}�^wo"����/`br�bY�j�j�$����~�-��KB��R���D̎��K유Q̋�[�bR�ǽ�������hMXʜ�YX�:&�Wk7lU �o����N��?�1q��ݬ]�%�R|A-���.k{ȉD�-�ɾ/N�
Ģn������at���-�vC���ЉF����Gg�"�i:��c�B�^��d�|ŪU¥�7N�@�K��s�C��uh���^TJ6�'Ѭ�R��`��r�!b�N?E�I���Tc��)��\&�x�$W1::���'�k��O"�8t�D�z1���u5䀱�Ų[���g�C�d�,�q��K���֒�x��)�R(%��O��v*������QAF�9���yed�h���ua�T4Z�^0�/uؖd�Meo"Ø/�q�Y[㠔��I:�樓M�Af�Br��\��׭�{�_@LrF�����0y�<ҥzdm3r�T�&V rh�5d�P����ӡ[1_��I-8����A9Afh����]�X�jN��f�SS�<3���!78��X���1Q��N�&��ByR��p&�*���%����~�#�Iv9 �X�8�FU~Nz]���,�OK��m*YQ�i�H��K/uZ�%chp�_�9�)���ðw� g��|Sg�a��7a��{۾Qg�݆��g�H�C�t���o�.�8{�Ҫb�rSZ��G��G��E�$kM�.��*���g131�׽l�rCkEt�"-YfR�Z��SC���H�q��e��鏱1�(�����K����ob�NjV�_�?�0���3��Z'��nf�9�@�Af��H�q�~@�+ڜ�4�VPzwq��u쀚�3@��R�?��8K�ܙ�X��}3;�\j��+r�����¬�
]/&�ҧ��Cm-ss�SA��v/�e2y�����f<Q��ك�}67�2c[yD�{Tb<s�$&g&�V�I�\�D�@����+eu�F"5d$paVx��&ϤY�JM��=�Jp\��v�s�Sq��	��YF/Q,F)dØ�@�������4m9Y{���E}��qC�D~�xM��Z˱� �� y"�R��}��r�f'�|�zq�p��e9|ˆ�f�0ʒ L�>�0�DbI�l��¡��5ߚt#!�Ž���0����_�Fzݐ�k����_��߅#��j���c����K�R��h"�W�fEϜA~�2�gr*4�tɐ�,��u�SISn'OD�w�̓�ϙ�YE����e��XDtCRØ\�Tl�%�dF�^	g�9�*pF6{8�(���"wu]��X�SJEF�r8&R��apBMA���']�rEѡ#�����wvf�1k)�/j�M�G��y=d_[2<�iJ"�k�ƕ%+Oii��^S�r�����l� v�r�,�FB�+�������7`PǄl3s.�GG�����|%Kl<�sӳawH��tJ2�+�Xu��P��gL�N�!��qI����KVa�o庒<ĉ������#8��cka�Ѩ���F,!�4�G~`)��~\-�⅟?���t���="������#;���u���s�T��T.,�k����i~���91F��J]3�`�b�3����+Ҩ˟|9	4���F�*�}�E���������n�l�3r�d_��EL��Ք@��y\9�6.N]E��۰��� ,F���lY�G�d�2Ӳ/�fu	�A�N��N_�(C��[�#���'#޾�^���?y�Z�Hm�ú[va�}w�3�l�B5�4c)$]Vy�q2�%�D�Rųⱃ���U=�q�Wo�����$�l�c�r�~�N�{� �PT�*[�w�B���L�"Z��\2��a04Y��C��ա� LTUԼ@�����R��S\b�U��=75���i���b��� |H�Z	4N;,v�\���йSpGy��R�r�N�'h��E�=��)�����}nfJ[Y�TZG'%�R֊�g�X�q�΄����`l�ެi��gU���Yw�;�l@��Q9�gi�/v��>&2J�D=򈑀f�C!+>�w�!��%q�$�Y�l��/�a���v[�:D�jͰ��F������mC:�^K�G<rTQ1�
��X;�N�P��_���̓�I��+��GϞ�3Zv�F8?����~(R'ի/��&b�	��uC:t��W���~UӮ�~{I�'�F�Ą�����ܺ	�m��D͠\�JӞ�z9{��A�^m�@�̬���$(,;��΂*��8ɴD�,q��(3�Kv.���[>k���� I��Eͪӓ�YY�P�q6K�PX(�8	K骨&�6�=�d��=U�Ҿ?;Ʈ�%��L�3���CĪ�fLMMK&�m4�%;���U#V��5,k��Ǒ��/PkCA0�@ˈ^(�Q�)&q�f��óHZ�:I4�$�v=�VC�A�e�w�%A�ѷ�FW:�m�u� ���8ƨd�~�b :�r�'�8yh�s���-�+��׶�u,�3[
q�A��ي���2�~�~ط܄�I/<�ǟ~{z���~�aH�׵����rV�*F�U�SD�j[���d�	���v��óޟ]���>*Ư��^�IC-��-u����Q�0ҷ���#��E����[c�l�(M��"'A�5V��o���?Cyf7�}�~��n��y�̯c!7
n4mV�Pf:�ҹP��apz��y,�z���bE~^�	�CJ�]��}��w`z7���}�-�\Gg�l���F��srt�����W��˰�6�Rec~S���)�_�G�߅����AK��,A�D�9�VE�����A�d�%I�b�<B��évv��Z&g�Mgә]�w�k)��t��\Eր#l2�I�Mn���4��<���`����n��VI ����+pR��mkBZFo�<�^�^ �Z�Q4�<�F�$xά�4��Ѯh&+
��t����u�$�=/�qE�9��b:���Җ�SĞ��Xͳ��U����6�O���ܪ�to10/I��sʿ�ָt�*�D���a��O�S҉��SF�m��XŨ��%���{rd�d��T���V0�9d����٬�q�p�bOx�s�%����q�]8t�0��N�Y
kzzQ��(5$���g#�G#�����1?�{�FWk�nX�NTg�D�앸����$yv�<�s(��(�� w�z�W�[~��,�T��d�}�vٰ���a��O��0㾂�X�*YmF2�Nq$jr ��2�!���y�l�����#���4G�*�V4Z��i��i����1�y�򕮵�Y��UK�BD��ƹM-�u'e����$K�4�����(T�]��=t�uS'�"���q|3^SJ�KW2�s�U��Ә�~t�WY���z��'P':Ն�`?��M�w7wu[B�N�hW::7=��|�$���/����9�2r�)Y��Xļ�_�+�=tq�lS�~�/��B����f�죆��k���d�ɨ�g��%��,��V<��a�� 
�|�A${:���;�g��*��}��G�F2��Vu�����Gh����KPT�[b%NK��ŕL&�ؓ�_Mq�����F�yY�}������G�H���$3y ւ���������4V���j1�]D��iL�E�J �/��(lY*_��=�w�,{��H:3��-������¨�WV>Ǯq�������/^���X�t �?� �KV�rH����x[��z_v@P��q�T�4�r���7arD��V�L>�$�lݫ�oc��J���Z(#�lK�g�֔���s����A�mK'�@叁e�|����Di�`������A�ڌLL")����1%�hnt\����.�Ǿu�V���8�A�Wf�q9C���&�*3ڦ����(9����3z~;8����0|wP�*�Y�L�3�e��P)�}�#'7g��s4��4����hZ���=�Y!�k���&�
���@������+�mF��8�FGN�|B�.��(��J'4�ab�ʪc�i-Y_���poy&�RvG�WI��03/v]��\��Sx��W019�{�|y	�Ͽw�/!ٲ1Z�4�C���{�����83{3:�����a������_�����n���W���/���g���M�P�}� 2� �m���P*f��ò��+�~�:���K�J�����)G5�0T�Z�B���'�<ɉ���@K�-c�N���dꩤd91�9���E��d)�Ǜ�.cv���(G�y�w(�H��x�&�'�y�TT�����k{��Q��3gN#�2#!�YZ�� {��ϟS�v�mY��Lm��T�=f�^�j���j�u5�𕣚�qU�8}U��`�غڔ�ƙ��&;WXd
�LN�U=��w/~����.��+�"%�KN���d�Yq`� �NyTc�.2c@����8�mFʚ�&$EKlހ~q:G����<�VKn����2;��?�����ɏ"�q9\1l^���� ;��\�,��U/Ⱦ,�A��q�+qTZ����e�8��3װk�	�z`QHŊ��g�BA�ʾZ���߁����/��n��»GJ&VCǊ�[u�+�c���hJ�RNű;�C?��O�7���b:]�����:t�Pf��2��6��.^�������͍�a����_�_���wa��;��zèG�i[.�9l߰1pαm2_���!8Xݶ�U���x�P��߳�V�%�ڹI1/�5+�L�bZ��E٫y�S���e?Xf	fv2�{�*X,�+�Q�Z�߼�����g�1�=�탃���vʽ�]�ؼ�˗��{����s��vM�9+u��*`s��g�&R�4�\~&/��:�����
~ay>ѐ��/K\Z(���f ��׋�8��~�d�)��f���a��%�����G��"�=Ak�LT�2i�H�Ց�@t*����F�a�VN�i]A����i0ȗ�%���x<�,�?P*��}�1`?�%���]��n���%�ȵ�M|F�z�X�}CX�t�}�9�:w[�����D��%L<!y����'�ۛ�"��.vЕ �	ߍ��a:_���D��9��o9��d���ٍ��T�|��C�^�
]=](Wʈt32�[�n����AC���-:� }���Q�["Rה�L<Q��
�ҩJ�pZ�X���U�_̃ɒ�fkr����!�%H����D��7���4�'�C�j��HH3K�d=�=J�윳�t�$�`����MD{<�������65>�JI�f�@&���2r�Uf�Y�,J�2g`T�
*�J�i�� ��r�X��Ԡ���\�E��n@C��U� AP>�	\�x��}[{�QV)hD�����UF� ڭ`ژځ�T�3��N=(���I���b��;�޺[7l�ˏ?�}?zw6\�z�CXz��Q��������� k��W0��>�� *_�=�Ч/��,5�̠lY�k�Ś<�Y�9��o���G�i�.��%KzW>���ht�g��.*��{�!ҠR�Qk����X�����Mת���`DVЖ��S�Z=[�*�CXy��̓L9lPYZn����lô1J]�V]y6$�tl��H�N�}Vq��8cS(ʵuoۊ��o5ٸm"��e�C!6��m���A�$�)�7g���GP�sp���c�#�>l�O2��V@�+kp���޻oah�*���v�,��F�#g.����j��0
l,7&>b���)�3ǘV�����b*/?���=�7,tmI*]���4>�Lb��u�e�n<3:�z,};*�b�ӌzY@����Z�~��G�~qB���u�L���P\���;�_<RTs�[�;3�\����R��uj����k��+	3f�5!6��/�Dw���9!���M�F��}���i�v�E�����~�	��{
�f��hV#�俏�m x��������o�3oHԗ�ƪ%�0r���9;	�}2��.��6Z�ӈ4}Z~��7������P�q)K]���W��������������ObZ��2�K!�~6��=��c��=s�4���{�=����بD4�i�fl߾/��<ZD�r���7n����%���c�P&
,��L�˗E��r=#a���T���9+��21�q�/� q��MH��2Q~�D4�q��2�o����.��)�̜x�:�X$���8��2mJY�&�P��Ē\��nq�ٌ8q9xD��U����4V��l�3}]�Z�3�-���6Δc��o:�ui�)�i0Dr��HQۙ���ӧq���q�-������ja=,m�~����T.��g���3�w�EG`�� ��jzQ^���%�E�%�4��!��6�K��=�#�_Q��][�v�8[����>��_�`�%F�d5H�!��� �U�W��Lxa�q���P��pڡ���+zq�7q��k�|t+v��2�c�%ݰR�!�z Rj������f���b$6� $F�c�}�������,��ō*�۷��eF��O5��鮵�b$F��Y�<�p�� ��Q͓fx��ţh\��R=�$uHu�Z1�%Cp��U<��@t}/�}p� ��#A�Ê����Oº6�k�Ř"U�Q#���-��֣���������~l��'�y�Qz� F�Wę�k��ύ�Xdj�%U�ҀÞL��;f�E�!����Z�=�K�G�TI_G��B�c��X�j�9qoI0���p�޽�x�4FΜ�`�{�v�Y���s��8���A~��b)+��f|3KO�ɪY��@QNQ��d	�%��ld���F���b|jR�kJC���,xX��On�V ��6���Z���q^+�B��̡\,Kp��k���?�ɾ8e]�U�=`�����AA�T���08�4|�h7�z�끀��R�B�#P��M�j^b�V,]��L�;�*��n�	�֭�����;w��Y�u��g�G���;K�H��	ZZf�5ܨ�ڡ�U��8��d�V��E���x<��l���+����ҋ�ѳn����������Λw�3��=�އ˗�����
	���j�*OHc��T��f�΃ê�����{�J]�J�`�7l*��$�(ϺD��^��j%Zf��Ct���P1����(���KgϪ��5q��׮E\���,��.L�a���IR�f<*f�ֿ�;R�xZr�I��\9���3C����u��̒9���B�e� �Dв�N�}ПC M���
2WX�ֲkd�C���5��9r?Q�£���#�q��At��$�gS6�?%җ�ͧ2�[ Σ�ҟ��s3S�0d����~��)K����~R�&!��z�0t�n<�݇}�m<�߾�_�~���0|�.L��:§�c�dd��d�NC	tJ����x���Ϛ�1�`�T�D�u����/��ҝ;0��\<v'���7����oF�m[`u�uo��r�|yVЦ7<��@�+��aO��v<��\c"���2�e�\C�ڐk_P��p*[��"C�]	��Y~uv����Aɟj������BM�c	t�F|�Y�LSU��h+��ɱ�����F�& ��7���A`D�'xv���!�y��Y8�z库��Y�"˛<�ko�����;\��|�!�֬�������`.��O>�\��OTE�̯���wM�b�ֳJ�ِ�nPk��$XI�{���KgB���J��iL�;�M��=���O=%��>��OᎻ����_�mm�Q�s�*�,Hf[CZ��V�����}312��ш��C���T��Z]�Q_.��>fӖ�[��#r�N>k!��03��t��:�W�]� �TL�c�媒8eĮ�2��8XG�C�P�W�E�A�lDi3<�����r=���ױ�ZK������>��Lru����<Y�(�6������ގ���sJ�=8ԏ��<E�U\=y
���n�*g!9O%/���>�s���XY�Q�s�nx��;�_��?�}H
G6���l�gݴ�{�����W�w���ɓ���z`	�x�U�d�^�N�6c�G�_��_�\/( ��7:<�z��F���ًJSA�eY#h&6�tn̾뤆�I�.�,�4��йw���D�J� �/,ȿ9��%3��O�3H˞zG�r�W8�J����\W��ɫ�5����5
�Ȧf-'련_qf	��H�ұ+���2���[p�^�M9�"���%�z�Q}gf�Z����Z�5:I�
e��گ�C��=���V��}M	���_���-��b�{�M�d}R��)���R��(�5��cK�\K=;R�X�c�r�a	|��Q�2B���Ɉ=Ն�Qy�b 㡄>7?� �y��_���7xM����7!%Nap|i��L�1|�!�����m����B
Z���*�7���צᦖ��*��@"#����[�p��?ǅ_��S3��K�i�6ϡ���3r`�DgM�p�@��\�Oi~.ePm"�@�==���i�����ŕ�����=ǤV�W��mźO~������%��ȵ���!�m�;Amʑ.{�A�eI`T��+�7{yo>��֭²�6Ò�����z�<�J�%���'LgU�9�q�IʬSD�k���r�
d��&�h�8YH	�l$*���sr�7����+��`�g?���a���zz
�voG��%��"�����1KJ)�'�A��ʥR "�'GFIaB*�"��ojI:��\2P��JB����ً���Dy���-���^��<�Y�v�mؼ}'N|O�5������F�,[���C�%��5(;k�&B� �F��y	@��sE�W�I|L�a�n:"+���PԒy2l���qڴU���UAM֕�-�tVq2��9y�ts*G��u�E���lV�d�̞j��Q�k5�0�3D���&`l'?�3k�7	�~ɹA�K� h|��L ����f��ZU=7l��d;Q�|�L�|?v�Z���~��^Gd�/����/�}�YY�������d_���縑_7�C狣S!9UO�x�O�i��B����6��=w�(B����m{�a�J>|�t
����s�8s�<��{A{�uqJ~$�O&���k	��V�j��L�cϗ�M��R�s��s�s 0���<�� �I�M�DiV~�@�rW��<P�A�b��3�RT,GYl���u�N@�X(��>�;�U2��咼oK�=TIK���������A�3'*�,��hyZ��1Y߀�P*p�3D�GlHd���NE����a Y�{�ca�y��X�r9��?G��U��$����;�,�6+��^�W�%fNT�3����1�pd㒵��<X��Z���5�4�S�@F��|FBՉ"Ν9��k�"�v9>��Gq��_����Vv�l�#Җ��v���36u��v�)���B)��}q�v�U�F�-�[�5[(cnbűk��G�S��-��k����N5�}RM�9���w푶��J1y|Q�!G�BW_|�K�Ѽ�C�w$�̲e+1/���h�y�8�A#���F��y���S	\�T	�"����mԎK�(�bd
�_~C�S���:~Z��}}�v��`��.����`{������b����Y�t�	�K�3�U,̼�&�$s���zk��H�����c��z�"N=�Ύ_U��M+лc.x	�R	}|.NM�o1��'lT]O�'�%�Qp�|�Zֹu�z����d��%��7�T��{n����j��nڽ'R	��ΥZQ���0'���/OZY���%h�B���Ak�2�]���=z������Q�^�L�}���ȴ���S%��f�z^h�4�wT(���X8����I���p��A!���*��.����[g��ٵ�#����~ ��`�)	EQ�͡����ڵ�I�C���5%I�nD�1OLNa�T���8>���p��{�=\~�-��U2@�~&q�ME~�j6/�V��QZVI	���;����p���'|�~�C��~��W;��gf���{r����?3؇Ub�f�<���p����s�M���0*��S�u���w$�4�� c$�H�܄ 1�����6�L<��h����� G?�gJ�8�c�Ӡ�7�B���+3�e��ϒ�r�N�V�RS���JN�fGSIg����/�zܰ�l�/E�<�M^�;Q�h˰��0F2��IpXe��Jii2� U�*�F�]�!'��(O���cT5e��5#��}�|�c�������#(O�ˆ��SS��Ê�O����OO�Πr4㊋1��z�M`�TQ�-���v@R. �Kα��0�,�|a�3�c��*гl���3HH�a�Uo ���C��u�T��?u�Y~�i=r��,�����ĥ�b��)y�u,����WE����{�wY:o �K�Z���cq�Q�Lo�  ��U���Qt��{��N,$-,{�Nl��6\���8��kpJ53�V�{ ^b�ڹ��/��k�݌u��!���i��g���&�س�����{�����pL-Lk��Z-�P�GG���P��3�h@�Y}������>'L+��:t��
�}�j�z�����nX�����������F����W1�a�����F�6��2S(#q���89q�*�
B��Ѣ�a�>�<��ꁇ�D#c��|�:�n�uh�������t�n�ЩBvN���ĸ�e@�T_��:a��9'�Qbcǀ'�b�i׀:C�|hġ���������e�a��!0�p�t�g�hw��F�vWUŤC�H�}'P�t�]#��z��X��
���&����Al:	��\$�&IP@$7m�(s�� >�U�H+-4e�������$��3Q��V�[�O~����0��;(��	c�o-t������k�f��F \.+�����ɍ�����p�|��eG�%3s]�'�^�b����z�Μ����˘~�e1����K���x��Gq|w޽��øx�*��e�9TШ�T��Vk��M�,H~S��ji�3�F�N�Hz��(XA�t�ɴ�� ������Y���XT�@Sb��a; �Ƶ��Enw΢�/�J$e-�U E4�*�ZS亙O��SYfT�/Bv���`K���N��l��_f֞�I�m���5s��l%U��F�fHD����/�W��k(�^�s?�>��A�峲�^q!ό���
�q0��M����,6��)�$ɑ;�-�����z�f�1%���Sn2NX����͉�X:[F��~��{IF�/`�B�RWp`�5��m:�4F����yy�w�4��ٌފ��L�ξW��O~.Yz;w����oA��a$����n��C�~T�c�ֶt�n�t�%%
����@����mz�:�/{�ft��o�(OT�oh��l���E�{@Y�����'Y~@��(��ɲ����fܗ��19�����Z8ޭ�t��kT$�*k��,�X-!i�3���n*�4��$�m�&5T�qy���3�9���]�
��r]�0r��DF�w'a!��Ό�����ć<ۢ��j)�g�9os�֌�C�9���%�g����6)j5�e0�J�^GB����cy��������v���~�j���t�Q�|����/oɾ�
XକPG����x|�>��c����7�w�$�
[��WQ ψ��ʘh�
@v�0���8�BP��u6r�:��[K�̾Y�o������ �S^�5�Q6L�U�n������9MG��$7�5���#A��`J�{�)�r��� ~tnZ���/}�Q,M�p�W�:{�yI�P+���N+�a�u&��<1���$��Gt����8����d��B��A:���t�C�t��#c�k���d����$K_҅�w��<���Ʒ���~�d����� ~��ϴTYcF����-#J�]�g��$�W��d�wp���/b)���P�n�ێ�G��aSB��L	��v�(	�\:�������I�)N��-�z�@Up�es�w]��Y�T�rǨH���PƷ�fs�����M������� �c,dh�#5i�(�]��7���s�����2z�ID�+��+To�#H*���%Fv�Jn�"R�<6�B�+�9�BE�/��,N�a�PS#Ti����O릏<��>?5��/�$A���|��q�
E$&f�U�"��F��X<b&�ڛȿ��_J��<��cv�a�z5�;�<[��Y�L�c�����A��eH���yja]su:�IQw��-����A�ٺ.��5Р�fY�Ь"�אL����a��q,��nZ��|��i�8|H	>(�N�q�VB���6�Q�F��
F�\	 +�\[����3��C/O��t�8� @��i�e/Ͻ��%=�HO�k)�-��<�e�@2�(�r}��s����4Zrm��� N+����>�ud`]�73kuz�-C�v+��N��;0t�-�<K8��AzuI0<�J����#����ћ��W��81qDdi����/����$���gi7\D=#�#�zN�����Ƀ8��+�~�.\�e�=rD[Qu�#�Ο;���n�m�o�AH�)�i�}k��3d����!�W=c;�$�|���q�D@9]��Q�
����TA<|�g�ry^[�~y>����1����T�wH��4�[֢μ��Y���-&ϖ/N����k`��
��x�j"���D�3`�{�D8[~�f@���U�y�C�ss�S�{w�ډ�_�����`k�w#�+�T�[�f���ǊAp)m����~��ơ��̬8��z�z�~]"��򝝷�ժ�O�͠0���#�Ӄ�b>��G�w��{<��
�ٲ~����<qE�<RYtg)�Z�^}C2 ��L437D��m����KT�"Z��x:~��-E�����C���dL˕Zv�@���(ѡS�E?0@�|���ݐ��� 5�N+����F�j���Q׀�R��n�;������<S��1��A��<W�(p�&�T/�f;MS�ϥ�x�S�ƎM��?�#.��ry&̘;�HD%�U�h�h�� ��0������nC^����@�^����f"�W�z-���ꅫH�|\�r���o�~y��$R�=h�s;��;���g��g�U�3�$2�Z�낫���3/��A��P������G��K�/]-�'0��S��]�Iv�D]��2It�8f���.z>;(���_�9�ܲ<��]l��&<����|�W����Q�f��K_Fn�Jy�up��6t�l3����|پє�0�3f���Kv�� ���]����_��d_���N��
bu`��]گe���F�F3E: W��v�.����'�>SOT��pX_1g�e/8 ~K���]9$�Ґ���u[��Ͼ�*ξ{X��"�t.��$��v&�d2	�� R�R�����^��k.anfA)~G��2<[ma����%1M�sg�T�rמ�0W�ǡ'Q�>��(�Z�LO#!o~B��X�+bY�.F���2#�.��$qQ*i��t�8i+�V��=hi/�g�V��U{��9ğp����0��՞w�[P;�����v@��8"dۏv�P|O�4�8�g�Qc:�n�{���}���Ţ$	��9r_�l��d:�vm~nF��8>����чF]��k����3g�W��F��\>�x���'4� ���:[�s*n��cj���@9�������?�-�DR3�f��S�x��Vu���w�b�9q�|�Z66mی�~�Q��O��_<��[�c��u��1O�O��47N��"F��p^�������Mc<	v	�M1�~���.2��z%a���6=\���4jn�"�K[Jn�l6��f�)���:?�q�q�f����ܠ��,�d�)|����g&h�p�R�����B�=��q��L� �ԫ��ˑY��x �~�!<����ȡ�0,�S�}�r���H�S%f"&��C5fa��`��jFyqns�B���d�o`�ug��`cW^�A�~=zO��Pg���~��+������S5��e�*�3-N�F~QQ�x�OPu�؆�J��8�8�faɜWu|l���x�=h��6���M*�:���T�`�"ٹ�;M�=C8����pv����&m�x�pa�8�&Y`l�r�p��(���݅�k��R�����C��7��s�Zb���Tf�>:��	r��@�~#��w,!ƳF�S�x��:�q��(�0�AU2u�,Ϟ�fqV�������b�#���[��aZErBl�E�H�#�(&��/k3q�$�}C���Ff�jY���Ez�)�>q��Y��5�[ځٔ�dH3�2A�&<8�"�o���+�XoN�{�S��	+���2�$�P��-�R	�d���k�J ��޻1[\��s�aM�@B�1$�j�*��j�L|�Re*yv�������y���5eou����!Ϝ�U���F�1j�Z}k'$���y�$�Y��6+I,���b�Fkg��z��r�4��D�Fy��I�*�G�P �#���+����n+i�~q��� �'$� ��ԕ�=&A��܍�<��c38��5,���AV-!�׾��~W>v�����[J<¿����~���r�|������ٹjbd%�pC�s2�J~��t�3���X>V8y	�S�ceO[7��|�.x�8��3X�a#�ߴU��K�N`v~ш��K��x#�({Q$d`I�ΏF�N���s���∉�$K��ܸA�+pN�L��oDhD�IV��X&���{*N��G��E�J����w�)0�򳵆#��F����v��缨cx����=��7�Y�!�d���6E�ٗQX�CoG��}7>���q��p���X"��ÊǓ� r�.%ƒ �+	��ɞ���}�c�&F�cIu�['d���J���q8-�X�P2��^?�W��g
��۱d�ZD^|Q���f[a���@��W��0�6����2����>���H�)2�%3��{�ǎa��1�8}Ӆ�:��XL����G�.����HgRص�f�
��2Vnh[�@p��)�R�Mu�Y�$�i�	(�6V��ǟ���A\>q^���߫ϻ<;�|"�B��g�~x9�U۶�G��'�W� *%������·3�"��(:&B�d�\ñ�\x�4��W	,"�`ٛN��b�<����K�LeK0K�tʁC���o<'������;aJ0d���x
�R�Ւ����p�4�^���@���/L��"�l��a��N$��qśǔ%�G�[R����~�c�$	�k�ƞ��`�|�� f�M��p$V�ɓŹI��i�!!�3+kҿgR���|�Ꮰ������#���uȽO8����q��r �L�X$�P�׆d��6�d?�8��� �ZD�[8бT�=��z�F@�l�p�_3$4�)ئ��IT{���Ȕ:S�w�7p�~@���r�y�a�sӦS�#�a��M�P*W���94c<ϴ� U�+� �C�j
1 fi�.j��*aKN���}����>��@����Y��v��(��HE#߬�����9���ZC�;����g���Ρ���?����?���8�(�XO�i�^MĒ�e�����9�X��c�PM���чp˞�������?��o���ӌBJ'^:w�d����?Ĺ݈�= �9p$C*S?�h�Q�������_�'�oi���ޢ�j=5eS�M�KƨP �a��=��]�H%�tN'����gy��o����ْC��m�s���l�_�ưB`�Z�s5����ő�U%�֪+NZ�®��?���<{'�=�!��^'��8��Lu[�d^d�l�#�hU�\�~���ʵK*�ù�Gf ��WԽ��k>-���W+"���;�ĻO��S��7T+��~��bH��Em/��G�4�R��?���R`�%��g�k��A�vN��ȳϠ�5�Ha`i72��I��p:��Is㳘�����/ Qm`U<-��<�:�mU�
��QBt#?�R/�]�����z��|FzV/�,3)�M~[/1�9.4}�c���cI(���єıwI �ypE�3[�E+q!�'fy9�����M�@�,�._��8�|GB��mhJ�F��\�ϟ�;9��e�R��{8���[>�����a3��}M��3��e0���)*��eIpܳT���i�H�#�5<��n	��iy��1�$ȱbI��9��ft� ABC>7��-N���b�\ˡ�_��T	�tV2��U'�n	�c��Z�sX24���1l^�_�����5���#H.FG6�J��jɨ��'M�Nq�t�|
r}Z�j�`�04�&ۆ>%��kQ�(9'��"Ϻg�M4{W���!��6U$��-����<����h'</(���x�n��&G�����
 �Z��MEѰiz���c�7��j�A���
��5��H*���Y����_�̧0���������o ]e���[���H,�=�Ko�D8H�ϊQ�My�����3������c#`�$-�;�,4�֓�ΞP���7��9��%q����z��q+�z���8����^�D9���g˘-�#��S�j����i���l6*�Y,�(Xj[k�`��Q����0Z"'���K�f,���[�K�x����ӣ�L?l���h���?�b�ى�%0�r� ȈF.p^A$�����8��F��j�@�J0�F�:.�z�Z�����0s�$*�.a���k���\��N0@�hY��PRT�V�܁=_|L�vcS�H�:�\��'!KIPRd%B� ��q�I2�JYq�k6��}m�N����)�2�jI<����B�j��\����~�n��{��R���M�Y	F�֬���;��3/tD���T����!�)I#:{��ڀ��iL�>��|���p2#b�t�+=4��b A��y���\���n��r,�g���&	u���B�H���;�^����K�9vS#��D�*͢�)m���X��ȵ% �n��l��ylܽ�僈gc�Q䣬XR���o�}��T�w�)J ����cE&��|Q��4�t�*�0�yF�2�6��YeR���-�}�?��tj$&�1�=�PoM?��"�oق���bD��9q�͘����xX�NN��m{4	�ly����`&�B��O�9l��V���:f�w���J��I���M�ɰ%��/_��O�B3�µ���[���������eYgd��v�@	Q�v���N⩊�zQ�Ӣ���+د*dnp��8yV�߰F��|�g��8�K r�y��*�i+pغ�-�R�ke��E)Y��1��ZA�^y�י���o/���_��-V��E�u;h���N��5�4�I�#κ֒`�u�6|����b+�<���u�T��_n6G{���4��Y .�ID��$�JEQ� �ͯ}`�W��?Q���8nd��!מ��ޏ�i;wyz�{��~ق3/��1q4C����;o��J�������WpA�pL6RRq�V�|��${��9kr(�r<,d��{Hux��}�Xm�	���҈v���a��t���8�nЫ6/E�߳�C��,A�'��\�^����i!}��-�0�U�^�y�� Kg欨c���t��2F@�Ք�6�%�b��%JU�j�x������먟;��#�0,F���a�W�5k�}���m�.��֛��c`���+�Ht�A�L��pT�]���?Kx/*A�)�5S�Go�=;����è�x&G�n�(�>-?��6y�Q�C[|ǻ��~]�ݔ=3�G"�3��%⚡�:��X�ླྀV��h�Ÿ7/>U����∝V�8��di�.�z��o�3�]}�=	X"�M�6Z�ȗ&��mX���/s�A��9�Ǖ�ކ��[��(�3�fR��-��Yjp�a� 4$����a�F�=��ܩ��K:>���hi�;�@�X
��	�;^_@E�~�14�3�;hE=ɽK!�R�%{�B'�7��bx�j�R.N< ��^�l+&α��5���3{f�+��2c��ʉ>ӓ%o�2��e0�B٫(�T���D�xd/�ZE��qqt�V����j�Tǜp�ƶa�#��g��d'F�,���>z/={ �����nD)uC�)�����rm�;�!�lX��װ����;_�*��w����W��?������ʵ͡�����9�M�xN�(Q��<��ٔ�Y�GB��=���ϑ�\3 T�����l6��z�A���vx���_'Fۣ��%l�=m�ێr�@ۼ-��6�Z��	�og$��3�n�Z��5ԉ��M�(T���૟~K�����|�m4�'�H��Y�1=4<��E��[IŦ}��]�K˞w�i��?��������:t���xY�5x<�n��N���v�u���sM6ו�#��ko+KѦ�~7�S�%3�������(+�����RK�Dw�#�|iD�X�r�.�&����V���)g��M4k�E����y�e��k31 ?(�#�d����	�9٤ԹU�:��8�i�fm�hD�%C:�h��ծ��.X�#f��:33�������}�����0z��N%1s�*-M�`�=�r�(���2��ډ�~3�N_��XgV���.��:����P��(e�|�����	���u��I�&�IK�bR�hXfQD�@v�6��/ۣTZ>?vZ|i�Bm�\3��,S�BL���<?|�|�Q\�xq�^.��x�[ԏ�=S!��b$kI�}��O˚���2#�Ϲ}�Ȟ4CdT�[g�m����	1�����܏�#hFS𦋸v���"J�0���^L�[���E˾J���������������GU�ODm%*Ҿ�8������$}9��k�
o� �\>�hO��shС .��&�����J`א�p�8�e�{p��?�w����w�2hTMvL���<K�fl�У���`��N���g�Igț��}OU�|um\���A�?s\�!�����(J��7jZ�b R-��0W���F�5J@�\-��Z���7��ۇQ���� V�1!Y����F�(������89=�R��G������*������#�K���ׯB'���*�D�*A���>_"ȉ�q��TY:o�����
��kE�U���R�m�&t�r+�8ݠ?n�{��+��@n~���cc��s&=���9�`��s�������k��C�@?hF�
;%�@�;��5G	���g�Z�ţ��>�_{�a�dm��b.�{a��	���s��?�zηZ�?E`�c�d�L'є��_�߿����v����?�ݯ�Sg Qr�_�]�ٟ�h�;]�����#���}k��~�Y��g/6l\���~:�w����"`)��P��.N'+4����Ѹ��:�Eį���m�_�R"���I{Z�:�m?k���./�3l���Lc	F�'g�igO�Z�pA7A&�3�
̨ۦ��z��#��Z��!e�Д�����W����]7�~�מ�	�����ˢ19��H	9М�e97dIf/�[��ѱ| ;>z?J�N�F.k	~b~A	+x�D�d�$�aד�+���5 �-)`9"�l;�G�,��w"/F�"��׌#��dl�LN�@��`�0h���v|O�m@sm��/�4])�_��>�a��0=?�|,��tI���O�;� �U>�%&ɂ劃vPb�X)c�U������JS��@��:��� AY|�V�~��k��|�({JB˅y4g���ݍ�@EV-�wj>bu����7������ċ=rϬ��}�T%�T	� �	����{l�3����i��g��i���/ݦq{�6�x�b�X��@�R�J�ڷ�����^������/"J��؍����H2+3�������ݑ!:o"�Ҥ��>�������_hMl�:e=����|����}���>�,�E-;�*]�%:�"� ���h�����6�j�Ɂz�W�q�C��mo�cgɛ��խ���rBжoѪxvz����w��n'etq�kn����<dFѰ4�U2G$���:��<��E�<��֬�nO
��Z�d��hϵ�%l?t@�,}���hq�<�XM�cA!z���\��Efp��W���	�lۊ���E�\���|\T�v�ڍ��<V���r�C���e�cF���\F�� �Cx���ը]}��q�BB�q�I�C�:O�:K¨H^(�c�Z�"Q��:E��;2�&RΆ��MDP�����e�K�:rK��DRo":�t���0wU�5D����G���=�y'�I@���׿��o=o}]4&"۪~�O��oǘ�l7��yY)r��I���1��	��o>�a|����H��X�;���u!�ݏ�Ý�������[3�>�����.�� ~�t?��F��c�c���:j�o��:S[�G���� ��P�8u���,q-G��4#7��N;y,�e.7��Dڪ�J�Իdn���`�c��ԢXc��wΗK5��=�ܟJ^1�3Ǫ�EVuC�-��V6"[U�[v������Hn����&�Fa���6n<�?�����ɭx���S�>�I�J���ô���W�x�\7LD�3��r���g�(^<s+�G� ���dF3���L����iP��We�(q�l�2����M%O�g2��O�"$Û���w6Tb�!��	�F��8u]!d�� �:]�2Rny�-(�݉���eU���8�)a�q��1�,��5�E1WB�@^W�J�`vy	�����^���Y�k����[>��^��%��D��}�{�������:OCC(Uh]{R��&�Q��4�m���
�疱R[¡�{1��{p���K:�7|d��hs,�au����C��η�Zm �����e"�8�ɱ=R�>@��#&>� �ڳs
��p��1v��y�v�0���՘��(��K�kЦ�����[Yg����s����b`�r=b����G�d�q:bt�"F����-�eV~c������Z��m��L�D�;	�N��I��S��Z"i��3O����R/��YCe���F��]�h��6\A9X#�n�9�o}죰��ƍo{~�GZ��|��E%L�ށ,�u�S|�s��eU�juE��J�W��2W��cQ�E>ZT teZ��,�Ӂޝ@+�E�Z,&H�"�~}}�kFI�N���>zQ+�NO�\�)}�"���*��>~&Ć�GD��d �z���<�t����o������|���g^����R�ť�N-?����P|8��t�#��С}�A�s�}��	���}O茟����������S����y�Yqr�e��bm�����Й�V,ڋO?�ӫ3���ᆻߌ�ql���>����HaV�<��<�Zm�tc�%]�ͦ�Qs��fP�e�
u'�$�um&hQ���v�!����~�l����5	�D$"�v�☄�;|C'R��U��;����s�����Kx�R)�tU�v�ސ��A2F�r�r���Ut�i��Կ���x�h�bk�(� �l�����<�r.�'�0njj��
.\���V;��S;�K<���sjr�����Yϑe�m�Olűg�%"8���^�)d��~��DF�������j(�LK�3��p�X��V�J����E�}�i�G r�wV��[�CǱ?fWױF$60T���-h�+"�[p�:�Nk��s��d�T�Զq7Wq��D�Ŭ���19o�(6V.�`)���O�F�b��>����tMZر}��	g�^"CKI��qz<7{�>V�c�b��{ތ5��׮a�āC���G��W�󵐓�v�]�%c����aM�bmm1]�r��RiDfe�<m���a���(c2t1Y�@T(����� �]��[c����jL��<�É8��Z�B�%�yV/�Q��G��JQ"�d�Y����3�
k�'���%2I�h���1�tc`|x㴮jU_
y=��Z~-�Dɾ"C1!2O�VK�Γ�O��@���chK��^�U��|D�A]:F<���t���t�_���<.\��;�� ~�=�Ʈ�����}N���v��5�0=����ĮhIX�g-^��t��2���u3�X�tπ�6%:M$�Є���Q�H�H@������]�f9�54�ҸJ�>5���Q����C��vPu�oq4 Q�.2��k5��Dt}��2�������| �w���SOa��)�?���<����_��x��ߦ}�I��'B���O���G?��wB����w�ۿ�3�9�<�x�Ίa��DgC;�-g"?��j�d�v��o���W���j��;���6�q�Ń��玣��0:4�}#�&�}���j�$���xC�Kϸ%�Je����!r7�7�"t&s��S��@5[�Eٮڐ���ɞ	���|"ti�
��95��TQ� P��2�~w=Q�C�E[)���XBk�#�bx�D��������đ�7c��S���|��K882�z�bGm�,��ٓ��q�f9��`!�2�ڎ��:�W�phS޷o/^q�\:G��Z�.�D �͈6�z�!��[�����<�]��A%u��Lt�;�i�`���}]�����
�TDF����(<��s��8�y��!R���1�s'N�<��A�����.�Y������[���D
�dl��s�sX�,Ʉ+n�ٹW��"v�xmб����6�t�C�Xِ:�[wbdl��N�P(�gw��xjL<$'S.��xծ���7��ZEm��pl+*��$"�[<�-#q��>K^�Gn�}�N������ �����	�/�)e�*�E��F[���e���qm�*�^���o��<��,�Z.����XJE{��;6-��Փp�?�!��p�����0���kB�CS�vc��.���y2,s2h�@^.m_��}2�Fv�aj�xh����7�[�%���a������kJ�o�<�U�y҅A��6�ssx�>�xy���سs;>������k�x9le���1,/.J���c1��|Z&S*��i;>5�J�U��Lx�ŵ�6�!��4��=p�i�N��&G���]"O�U���VŊV5����âF�L�/*�K9,���i�NzN����߹b;�X}����o���o]}�kX}�9,>��t!8�!,͎��I�9~�u�ƶ��!K=W�h�T�!sC�}��_�0~�����*�KaB��l���Y��5_.���ƿ���Fv��֥?�".c�]w��+cr���Ƕ��/?"y�R~7v�؃��$.L_��ڊT�7�Uz��$�����~�Jbj�Z��i���]���|[��#=X% /Tވ�����Z��%�u�:��cO�{Q�*\�`E�<yl.�3�/����5w�]w����?��x��_�W��Fڜ�ZY�e�,����9ϝHf�w,���/�Q�S@d�� O~(�����!�%_Ρ�"���M�2j��C���:&��`�������I�����]V�Z�������6\ȰO{��'���~�XJO��٢/��\q�g���n&/�*�Aa�N�}�.��A����qk�]%Jy�L�W�U1m�6�mغm'���͞�ja��Q	�&ܖH��<��U����T�{�i�BMV�k�QW�}E�b�qH5K���7f�Z{���<g����� ����ym)R�BJ�n�Bs���Z�<�
�F�`emCt�3,%*QoG�l�nAϐ��m��Mbb}����TS�
�P2���OЫyX)�t�����#Okm��ntr,�!G����4����F�m��F5Z���!d���8���d�]s��ULn�$�d;�<�J,��9�V���y����;Mx"� �	���u-I=�a��&J�,V�:����auq�z���?�><������n�i=��@׮R� �v�����[2!1�St22Ur�:����jS��$T�����WK�-dx����Լ��`�ݍ��A�x��%E�\)�מ��ص�A���j8P;�+Dk�\��z���q��1ԯ^���E��EDW��0���z��h7�b�)Z+�ފ�o��Ja��[{��k./�ʯ���w����_��k�	��<�*�|��Y�#�I��Z'��T�r��2�t��bep�X����ڐG�/a��;���އ����'��SO��'pp�M�������̢�^�:��VҔ�l��!��uu���XzZ[Z�r���y>r�	�ی"=Kp��HT;��k�jִ�M"ؖ
�el5��@r��s�*mt���M�8��}D@oz���ʛn�ܷ�᫟�2�����"6rD E��2�l��V�?��䩄��nVB~���=�t���!o��6JX%r+������h����D�������h���R�D�\�ǭSI��%]Y����'����!~�_f�J[K�v�C?��x�|�{&�;���Q��t��om&��s蒇B�g̟���mي��u�e�rY �S"�Z�r��
���1�}'*'+�U�deɳc�Kꑄ�#���CW��pA�tG�O�&�h�ZJX�!�<[�� �{�QW�6+�C�5��9W�汃�E�px>vM��b�d�q�Ȁ��%zz�����	� ������ƚ��KE��%$d0i��xUf	�r�i�:T�X��oW�HF�W��Ed�"��K��E8-�+�X^]�u��9Gx��

d(՚K(!�-�|4�3��PN��=�N�vS;w�$��ҦD`y2��RK�u:�MQ%�y�|�2�\��Z	,|����n���YQ2����:榧񊷽o��.��f<��3x��%�jȃcF�*r3	��t�6dD��U����d�{����XO��A���d�x!f[�0��]��6�Ox�F����K�g��I�y�^�'ܢ*�?\`Ƣ.(��E�y�uN���Sx�=���ފr���������`��9��K<�����L��}8������ȱ�vv����r�Y?��A��_��<�����FL^h�)��)R��F܉��������ՙ��w���ӽ�1��������}�}���Cؿc>�/|�k8�2�lߏ�S�02\�z}�����;\��jK؝7PU�k��nkB瑚>��hq�XW��-&���Q��Swǖ�v)v�,ݒ���X��Dx�[n�'O��R��rm^1W��&��i������[^�W��0��:�~�S���S�u0N�í50�pn�����rې>�t�3k8s����g?�I�h�Z����S�:�,�N��|�D^z$�L����sΒ�h��_Ԯt����qk��6�y:�le~=zn���9�.;���`��f����/u�p�{����l:ol	q�-t �)�h���!¶DA�cxf3�u�r��%@YT�_�����o,$�b��U��WՖ�{G���s2���Gr�2W�-�H��$�+�U4�[.���1I�%��1�c+�A�����:!��k,�)��f����d��ɵZ����Ȩ`Տ|TYÝ�Z)�$ժ5�7ZZ�͖�1BNR̙\����ݤq/��똫�Y����B6O筎���𑛰Di=n�Ѷ��:�e��|Aj&��d��t�8��ٴ��_\�Q�9���Ҝ����x<*��bA�L'�*{1�m5z�-]	?�n�2�~�|��%<�ǟ��/�u?���C?�.���4�x��x����ؘ��zV�G�pQ��b}mM���X9OD�$������<U�W]���'�.I�z)�4�!�*����:;.F0{��tt�N@�t`y�1�YZ�<L�e����;���݇Cd��p'�xgN#����O�tp�oQ�=90���DI�b츝��RtM2y4ɘ���c������܇>�_���@�,��P	A-A�I��Zx�m3�-C3זW��5�ݕ��7f�t�N^]���a�=w�>�Do>�J<��sx�;'�}�ǂsz��ynlT�Vis���N$ϹtKk��:�ձB!�8M5�n���-���+�nu=�$vt��rsd�� �����_j3�L��;(�Ja�j�.8;�m����w�+�y��o����D������\���^t�כ�yg�mϑϣ�S�+����C�%%b�75t�� ��D7齧����sW0Y*�02+[y���Y���7d���Y���.@Qz����Ԛ_�7��I�lPߐ^p��p+�ck��W�!��6�.�CmҪ��sDNd��>��U@&F��ِ��%��Ƒ��sG�3ޠ=�H��S(�H�=�[�D�G�r.�'C$h6epL�Ɋ�~��[�2��p���[��)�jx���	HX�F$G玷������xEW.�����6��&�=��";&8"_�·ۤץ���i��!a���ÎH.��t:^R��'t~�^%/�.�s@�T�Kl���U%2�F��KմW�3��s��Q����:������*�^A"C���$��َJ��e2��Qʉ��C?Jd rU�<H�m!-�;2P�f�9{����WO_<�T��x�����daÅ���P��qk\b�H��$� o>��Y��s���{e�Dc����ǃg�1~�0�x���矿�ϟ��Ǐ��ɓ<�[������l�kѵ㱴��bh鼵�Hw�:B��l�
����*����fX��U9 V�
IT�C"Z\�)Y<z����4[&�{�[���r��7�oz�L��Ak�o<���']�G�N����7Z5g��X6���j��[t�����œu�3�k>@?�k3d�r0��7�?����|��-ϔ�,aA^k�H��t+��#�]o|�B����߾�����6/�c��CXy�8�n{F�o��5x������8�46�e�A��stb#[ƥ-��h���b��H�>y.2���t�s��}qu8��r2W���@|c��{D�%���ƺ���B]D#���y�YsN:�� ��t[�o�=7߅��|��|���<�-\�ַо|#��Y���jn�Ԉ��fe�H(_� ����-/�y����2��"��Wfq��\��������8s�8�2�̎�p7y*Ǐ>�m���1��w�A�ɐ�E��6�8��ث5p����9�@Ɔ�:,�K
��_�C�_��l�^�7@�(2O٣��q�uvEHe�����U��p׮mB�s3���a�J���I3��p����5Ia��$웣�;$�^�6�O$�a��hUμ$X|�$&ￇ<o52�z򛸋��w��_~H" ,V2H_�_~�Gɛ���w�sK3x����B$Xj�:���>7�"�y`}{&�N���\	�C��wȤ����Kg1�uJ���W�k�N1~�*k�̉p������\!rj����c��v����:<���=�0&qJ&�B��..��ZJ�H"=ܚF�h��6oD�k���k��q�/��}܇�F�<�62EՕU4��v�ӡ�Т��6>	��>�[2�ط��q:���ψ�[��x�f&
e$k�-���ID^�8�n��S-��w�LԷu�>L�߉��f�]����J�@4����2V×O���+��{��8z� ��i�:s���2��[7����@�Ѩ����jH�I�G���O�ӵ:\ڞƆ:��S{��'SQ!��ܜT�GZ2�Ui*:n^�Sdi��D�\'��Y�cC8r���կ����ڿ���`�̋֖`��(�\�S��6Ȣu܋�����I��~_,;�;t�;��B��xh��_��O���a��������ԏ���"��"�j����t����e~��g�����f��2��e���Qd7�����C���qL��jL��j���𺻏���x���i3\�}͒g�dB��1��<��Q��<�Z[-�P,�O��x@�j�
%�ȹ2��c���v2Vy
��rQ��2��s�9/�3�yn9[���;����ކ{�w�E{q��N<�,�9[�a�n�a�y�k밫�I�IS����U����]/�Ms|l�/.�P��{P��������(n������.�:A�ٰ����{_\[���v���\�
y �A�j�a�%:��ʱ�l;���g����7�����L�4Ʈr��B,���G!;P������Փ����.\�ks��I�$B�"��(A��d�@������kצq�M7�};�`y˳�&2K�r�*��(��[$c/�yNP�C_:sS�U�#��l��h?���p罯�։a<���brκAk��������j7q�8��� ��"�WN_T���e9�A�G�y�KdH̞z��>��7k��x�I�G���C���	1�Z�5T��ɛz�[�@�6p��P&o���
����	x�P<^׶�Z�.z~��@_[_
1�ؘ�\����}S����kg��Z)���X� �����.=�B��=;&��Ï�Z'e��Fkgai^z��t�k1�sp�k_�0����pz��*	����KŎ�}��.�j�t��Y�⦛��"X�Ci��Z#�z��і��Y�����k3��ԟ|�>�E���7a׫��-o{;��><��i|��Q\!��E$��r<Z�21�U[����K�C�J�F�A:��D������NiJ�����?7�K���~���{�嘙`�S5��%��Zză��ȣ�31�L$pD׃��m��Y7lɊ�]:�7A`�O݄��Y�(�÷3��0���9��/V"��UN�d^4D����ؓ/��r���F�!?���$�^����`�=ԡj�\-x˪�M��U<�b�?S1j���H�o��p�o��I�4��7��E��g� ��a{f���v@���-�	�C��{ݢ4�1Q>�����"���Y��n9��ag`�&D��F?�5��6����_G���:t��4�MI�?V�ar/C��� {��ʛ���RCƍdi����f�_�Qf?�Wf�>��U�O��gcc��+-~w�#�������%W��0�_Y,��9c��)"���l}�L�@^N��w�:gX8��R���M��� ��g��P������7:l)C�>t�� /d�5v�^N�x�L����'�Ջ3�z����j�wAS���c�f������gg��lP&��HV8�o�K�mP�������O����=���MB'J�>�t��u��mk$N�ǯ{܁h��D�@�9���?'�z��E�I��/&��9l����툙98P�N��jԯ�_Z���=�*^,���C'ʨRzA�8������3Ϗ`s�*���&&Y�o�Cc�t�tV�K�?�|=��Ƭ~���";��`\�M��`4[G*[��h�2�rs��-ƨ�ᬇ:/�����萤��F����/>�u��_�yK�		�\a�T����hzqBG{TŢ��_��_)���f}��xlC���C�9Bi��6�b�sPBE?O|Po���я����.g��M���i��.=��xS1�g�^��Z�R��g�=|�����w��G{=A2욨Tt��A���Oǌ��^����Y9}H���3��ȷ`nuƈ���U>��W��[-�O���dyA׬'7�BG�;5m4}������:��^�-�2���z��(�Ka:c��f�f�s9���"���ԆQV.�W"֝��J���s�����+�2(�Ћv����m�9-�
jxC��������ȅ& ��`j��N4���`,��7�R5<��$��3u̿8c"��(TM�A�d�it]g�����5�Тp�m�\5��쿮L|��v�t�tY9r��Q��@��c�S���D [�^z����s��M1�xK�i�9��r�n���>�Y e� u�T��v������@��s�$�e\D��d������ C�l�M��H?�)Ҿߒ�Z�v�VI��d��ͻ�qۓ��7�i�r{&�V���������Sa�s~��=)
��H�3��FR�v+��M�(-n�lgM!�~r��h,�68�f����y3j�?��u�&�\ӋlS��Q�&�@4t����E3z7-�ߍA��~ouя�!m|�<vPb 2��8�5�m�T[�[yd�I�2p�<���������=���&/�q^�(�rQ��#��ß�'0ҠHF��Yс��Hь75��o�"��3���@���Q�`�Ǉcv>iBv^X������l��X�4E ׿1��K��H�@А��TD��� )���� �2d�V�d�h��zl�$��0���n�QmR6{'�N�`���	u7�,ܐN���Co��}Y7�8J��/���f���)P�a8�g��꿘���.|���(%s��$�U;�w��<���`J�
 cqgV�%�+N�9t���Km�[]╵s\D�"^t0���GX��z�۵�݊I<���v&��_*ro�z#�Ͳ��iX��,����\S$����:ĵs�Isss�Od���M)]��)��7���Wn�����f��m�&�Pv6��"*d�Y�j��7&��K���#��?D�T��_Ѣ��_�>��?�C���t<��e��M�C\���o1e����y����h�����f�Q$n�wf�6�i��zԾ-$c�ۅ����t�bWW��I(�ox�=�fȺ߭9�F��ʜ2�~Ӕ�sMˑ���0_��`�`�� �T���b�w�@u����J�pdi�O�j�����@�ς�b�Ҙ�+,�_g�u/c �Nkz��*_:b�~bCw#Y���_nJ$zy#	L�}��$wv�7�Oc� xPdBC���J19�|����b�$�^�¬�\v(��$���m��?t)P���;xc��x9+��(HD]�lR�m��9��Y��:/��@��_k�u2�}?�.7Z!��E�
�t�������7>�s� ��)��3��+����q�g0�bO��%2��\#��x[#��Q5ʈ5m�[2���x���-I��,�S��뫻i�e��i?O������Q��p?�(�F4v�� ʝ�E"�m�.phP_(3�N^�����E�:\)�g�d��b�V�K<�^�S~��ZW�߬>_⧎L#<d@z�CK���p��M����ΟW�Q�n�la*����d}=��4��J�_3N�w�߾H+�`��@�H�|��.V�3?�"��3��` D5�$��aOtN]Ǫ�6���xx"{��g�4�fʌh�#l��+M�W!:�V����=gۊ^v��ԁN-l	��5&%�-�ןr��7<F�s���I�tuL>OD�]�f����aU��-��
g����H�
$M���$nm��)�����#�T�:�x'��ZMl�)u�0���D�ݐ��IYs ?h�zxٓ���b&�Ǵ/����*�P����FԻ�?1�=X⫚0�:��|$����C��C�qS�e���m>��.��*Zr�k7��3�����L���j�0��s=�m~���4�[��ŏ����~lbr=��Y�{�>C���N�ټ����ޛ�T5�}�H�8���Ep*8����S���l��i�2�ٮ��_�^�9�N���K^���og7R����^��W���^n	�A��Kv����	�<�����Y��y��5���/{�ٮ=s���Ż���ZrmU��A@��O����TxҀ�&ӟ}^8R�Ar�����o��A��_"3�%��W�<c+:�ѹ�Ʈ���SV� �9��Zin��kޡ�v�~7m!��7��8l����T.�ii�j�g|�ͱ! �q=LJ�n�_�9Pt �K5�C��ip^�p����}��ݏ�>�]L :لh�A�ܞ�'��ݦt��ռ%+G\��=��h�j�:d�
Ϊ��A�A�Glh�8T
��!տ���u=K�m� �ֹ�q��,Jk�hO�/܏$�h���St�p"�Ѫ;���8�u`KϚZ"ؾ��eV�D�Ju��؛�2��Q��s��̙ό��6�:��Wi�����v깓t�� I<�?��j�8�:���K�j�������?��F&%�Mk.�5�����uY�xJ �1��w�����������Ů�&���aQk&[@��OO>OM֙Op�ZqT���Y�p$F����M͢��	q�I�[���Q�F,�BIS�~���v�/Nps��������|����l&l���)j �-.���V�ZNx�R���N���:g�p�/�B�v]A��)V�C�{n��~9����'8��|�,B>yc����?{�y�\����{Uy��Y9|�_���i�[�h�
������+�r�Ƌ)��������L-��{�"ȱ��H�ƕ�ss\]�@¶���{e�{������d��G���(�� ��X�[��p��^UF��Ww��ɚ;����Z�3��^OG)�d�VZO֢�rExz����=E8�ދh��3r���y]�nԿ �V,)����5tV"����}���l��{���E�o�M�\[�$*�>/�dv���w�WXI��O��S���&���(N�v��u���"����ʔsO����d���]�jf;�"!�/0�?���;�7���͗�7��h��=E���<3B�L;p�G���e�h��לA�{�b����W���}��8Ip���*�~�ס��3sO�vi���UN.������;��m4�1ګ)`Eh�8~L)�x����V��h���~��{�-�'S����'���m�a��)t����՟Z-0�}��?�}W�K���ohV-���>#��P{���ƶ������gQ���_ژc�W��"\m�K�����G56~�P�IL[���:JR�c��%7��@U*��Z9Ŝ.��5Χ�����tT�1�u�rNK����<���'�j�8-p p���2�&_�&���FN%�ɂC�ϸ�JY� %��2��b�o��U��r��5�]5ߦ,����ہ>�&eH�}��+��з]�w��o{�ˇ��/�����=�`M}'� �H7���|z�r�mRۦm����D��>�H�|}|�4���*��q�g�]{�]&�wį켐�(�("����X,��,�k��^H4�aI���B	U��Xs�����c�ϫ����^n	P����JE�hy����kG�u�Uъ���O����P��O�$� -��ȧ4�W�Nd�Y��KC�Ŧ�ΒI�ky�\�Ž�g��l��~�5dm�ɛv�Ѫ�>.π�_�q��V�|�n�Lrj�$�М̾�x���e�x�-��ǟ`��[�E������gFྜྷ*����(�8{��|K��f�]�u�]k�j�a#��b��GT@�Ԃ�`3�X�Ee�,k��\�@�Wm=Bt���-�ո\����gb�M=ɐ۸G8[���m��Nڀz���x�o��(�j~/�N�]{\���*�d��z�)�Tf�h�O��[bΣ�PyB������=<��]x��_�߽�ʉ��>Fq�s�2�U�����bF׶�!���t>��{w-f�ԲcT���D��Qan�`���ҜQ��wǀi��NgY�;����f�1˥4k<�X�n
���>�msu\�ӭ�5��l�	�yP=�O��s���љ�b'�'���梧*q?*���Պ*����r[�����8Kʵ��~S;�5��2l��-��eA��DEhtG�����'��K�v}����B�3>U���b����NݮE�sA�i��t#1�P�8�I��?s?)*K���\�9f���ce߃��Ȥ?�q��T���W[��(1�W�L����_z!5+�/���� �#G݌3�����Ѩ��X.�_k��$~�(�EK��܃��&����k�2x��<#Ӥ��*\��FPb�/�& �e-�[5�_+z�Z�k��s�&��2�C��y�#3���ӂ����2Kw*��BW�!P�OnJ�V�U��p�V�H��4'��Y10�k���^a3PI]���7jD���%9V=H6p��r�/XdZ�V��a�9�uw���A�1��d�|T�0I�@,�Q�"��"-HI��RƖ׿��~�v嘜�p\%"�]�q�J�96��W@�F��
��Y�#��~7�|�����)挰�
,jc�:����fQ�`lvn���Cv��03�����丂�%�"!W��/\��^�y���
X(biX譳M����D�d�����Glc��
�6�,B2uM�u�݌xJ��o��T���\j�g�v�R9�����7� ����߾�o�OAzl�"��]�&N�����n2z"��V��8K����q7���W��W[��OOb�Z�2���q��8FR+�BG��?*�]/��E��S�[�tI��%N���u��P��`�6�����j��%��H��[������GUr�ӠUU�4�k�s:����4�X���Ѧ�FlI�Js{�Q�	��ᥗN�$�������J��tb|vj�<������;uh���u_����+i�Ѡ�z�xr���w��N���X�Ĵ�4�P���l��� 6S�Q��zD:�Y`[wf�vE���4�e=��1�Զ��#\W��^Z*��ʐr���4��m`���cpj� �L�Ӻ8&��N�<"�Ajo�ti��xuu�����E�C�em<�%��B��-HpYzƍ��k��Z�\_������Ed���㝴4�@AT[H�C�a���;\,
Y�Rh�N���NqK��U�f%�*��@��u�(H�UKA[h�%����W�b��)~���8��p!ŜK�C�XU�b�8��*�Ȏ-SlKW���@��F.̉?~y���>5���d0��+ʳR�*۾me��su�.|^�C�f��;͉�e���/ǔ8i���Q$�$! o�����>@��i#^��$�*��������#��®��ա
�#��83E.�C������CN�??$��M��q9������� [���h��4�*��Ns�:�>�1�[�'��+3�8�ٰ��w;sI^�D'�t�-�zD�=�1{n��q��)G�re؆i:�ﴂ�d'��(M���Ɔ�-]�ғ�4�T&:�TZ��rB�$T��R��������K�rQ�]������e�F���'k�R2F��+�0A<���f̌����-����J�I���p��=��"<����Bɫ����⪰�rv���L'C��m2W�k�Vr���������ꓲ#Q��O��75i�X	���&�᠉�zҥ�D�	XR��)�8<LL�-��m:)h���������������7��W?Yą	VY�ĂO���[wB�m�H���" ">����������|��B$����K'1{�~��C9J��D	 Y ���i$H��N�S��/�>a�%Q�K���6�����
&mʜ�=Q�pW2z|�n_^,!��JȞh&NI��Sq�f��qχ86�ݨ(����"���U�Z�~��!�G���%�����4��E�,f�>������e�hL������1�I�_#��C>Yo�(�����N��(֘(/�X{�C��%�*)d�[j�y�%��,�8��H��?���xG��&24F�]x\�M��ry��R�Aq3-�YR[ӯȘ=w<��w�8���'A���.�ˈY�_�9�^�;�MB��=��S�}�f��:���]	jI�\�iv9nT~�VL�p�����ҡ��>|&�g{�J�y�ԕ���������A.�*�P�.ӕ�d��H�4L���O�ҶxK���|Ôsd�c|aKit>4��S�1˕�ԓA����Y�CW�c��?��F�*��ef\> 7�7��hOY&�f��\>��H��6�`@��a���c�R������D� ��4��T$��a���Q��H�3�V�������J��t�m�'��cD���?���bY�X�P�xq����al�`�5�����{�G�d�'��_9\�Bt*� �|#Dxe���	9�m��Uf����_^k��;�j	pN#��ayj[a����&,��R�l�d�Y����g)N�꒯s|>����˗�x��Nj��>�?���~I򅔪��AI�3�3\W��J��O��"9�?�
�WO�v��P�ޱ?_�00�f�g�"���ͣ_�c�|V�{�C���62�'������=�E�q,~��~�Qy�BI�G 7O[ܝې��O���U��R�BNU�HS�u8�YF��*��E9�:_x��(A�MWs&;4
.��2�	z�!}~��}��ܳZzyx{���k�׭����k�r�̽��St�LW�v�m�X���$�tWl��}_b���4�أC��dވ��;|�6�ߑ,
�`w2�a
Sa�æ雑��W&�R���H�h�E<�C�D2
��P�]V]���/=�X��d�:���T��+{���H|��xM	��~ലid"��r�qV7����qL]�a���'��o+J�f��;�
�Fy[�{�٠��v�^��*��6��M�m�k�Z���$*L�7������?�[K����4��~KHz�����l��st�z��-'���c��UPl.L��O�@�<>�4S�Y��7�V��mH̆������E�~Q�7h�8�ӭ��0�ES_Ro}i�y^����%��1���CE{V���.QLK+�E�����S�5�
�� +�̃�GdX�:r�}o�Q�!1��:9����\�+��Py��������̂�C�p9���ۉh��Ӑ�'K=��׳[��͊���hs�t�PWO�ik�=b��޲��A�'c��*}S���ZY�UPe�@|�$�xu>���.��2��B��`T���&�c�׸X�G�^F;b&��?�,q�}��O�	�����d������M��k����=��hg"s�XE�������ΡK{忴(U��2��Y,e/�IU��(9�é�������o�`�b�F�t�	µ/�#��b�� /��Ч6c�1c��ht�mZ(@�}'��D��u螝3�:v���C��zo�U�܎g]7BJN.p�T�4��p���m*�O��i����[��H+F��V]�X���m�h��XbD��R��(|ix��+8��
y��e��5�ĝ���t���pT��J��R�'� �6	�xA��5����1O�wo��C�(S>�<|�}�<�;eM��@Y�3u�s�(�� �l�̈��Oz��3�jd�QQ�>�	߅�,P��1��k751�ޚ#O��&t/^"�� ����4U�G`a/����B-Xˤ[�v���!�q��U�C�&c��ސ^W�@���D���_�A���h���8N[��h�T��˼؄蠈=\�<RO��8|N��n:|�Y��C���lE�*w`$#6�a� �.d�tZ�)�5,�gCauu)�r
-�����mj��ri��<"�&f�iۙ�kZr����g��O�R<�a��A��/v�O_�c�H�,�Va(�%����
�bB��#����AS>&�\ٹL#����Y0QLLC� �M��\�uC��N�5�C�ݎ��U:��U�s�j���UK��K�G[{v݃��{�}�2���	��.M��]��,.���q\I�3�.K>Bh蛲#����9Gt���꘷�Ԝ*��
���wc�zڕU��PE}��Yf��Q���w�ݸΐ+�/�m|DT�a�"�^+C�f.-#��g��pSk޿�q����0�R���7��%X� ���<�0/o���^���-�l�B����_9�h����	(b˚Êe7P�޻٥����A����Ri�Sr��b�U����f�,�g־�S�ؽ��X���`B����l�{�GF*�[�&����OS��	�u�剢��t��}W����d����N�z�������OC+�b�Z��tJ�*?G>6�wOFN�SG��Y����߷�T6v��B;����n��U��4�Y��7U'��J�.�#UR�Ix9�л�v&>ۂA	?8��l�}N�_-!䀲qo:]xX��z���}��G�:|�_T|u~~�})DM��*�V
�R�hR%"�e;e�ya�ֶ��Z�2�Y�_�jEۊ��
I����t�-y$I�N칫���U�9�7;��<���[[�z��X���~���'w�I7m����W�ZɢU^���͎���< �'�9��/\U�+;��g)N����5"N���	��)�.���1�򈏠9I��`���$��!�cv�7��WQ��1�V-y֥Vg�U�{WʓŜ�m�$r�fe5uߕD�3�j�*? a<sT%pi����]������ XIH>`X�>TT�͙.�b�Y�0�oI�����U �r��q�u��^�� ̧���X����J�S�K�f�X@6w���$_�
R^��$�9FO)��i�7}ό�R��eX;�S�oĉL�lL���z��tI4*wb���^�5������"8	2������&Һ@`3���9��4{�}kU�p�o3�plM�gE��� W(������JP��~ŏ��>�T ӫ���r����O!�Ar�A.e`��+]�O��s>)%����$ǩ���(�"�x(��-�G��=�5�j�&�.�6`�$�x4'�kd�\��maqV�Y�\���4�������VMtI���L᯾����Ӑ>	cR�7渷���M�$Sߧ�D�ԑ+Z.�� Ъ�UE#�Ъ�@m���'[�#�a�B{]Vi��L�7�he/�8��o{qԚb,+mհDk�k	�]�J�Fq7�����텡�"\L�c�2�JV�b8�].{j��@��9�z#_�ƾx�qx>����W���Vo�]�ԣ�A�uw=Ɯ�S�L���0���k֚*��Ż#s|��˖���Z�zv��V��k��!q>C�@�f(��u�ַ4��MK {Ռ�l!Qyg/�ڂ� +�Z��
?y��oޏvM�R�U��^ٜ)�Td�1]y��2}�(�D������DaH��G�� :�Ӟ��eb���y`���b�qgB���`!�&;矍F�S�W孊�8:;�C"�hY��XkBA��.&+��m `��J�])N��OÊF��a&�LbKcx�;�AS��Ju���19ލ����X+V��d�Q'W�_-6�=�>c�{�4O�w�ӽ{���߻6��!f��?�<Q�>���V�\ �
9�6汿��>Ș?z%���`r�M��Q�B��='Kx��'�4}]Q�X� �{���4-��Oh���2��"5�ؿr ����=�ꂖ
b�G�kq,o7
%6f� )��o�]3��==p��w�M�_4J(f�Դ�ku��	Q��k�ti��������.�����W���/�`���}*aR�E�zg�)����cJ^x�,�z�e,�60�j�3R�>{8���,;{Y����O/j ��O#,ұ����/K]�}q�Q~$O�щv�%�;��*5�['_�8C�����w� ��8k�T@���;�|���nz�:]o!A��Oi�鏪�ѥ���y�+P���v���%���44*%4^M���קS{�;�?��ր��pn�}�b�YJ:�N�:��gl>_S�^Ó�Yy����k�X`��sj��Ւ��x��P�k��i-�S���:�溞�s�\M�Eoy�Kj��^ph�����}R
�ߐ��y�Ɠ��bSڣ���=?�a�AB7g܉ >��MdI_�P@N���fY2��񭕩M��3��v���9�k���RdHi[���:;\ t�d撉Bo�{�;jK���E*���Q|%c O��Q�I:?�|P�t���H.�o]�),b��Y����Q-�X���o�c �е�~�r+_$�3vN�b��k��=~����~��yw�y�Θ�� t�*�����/y�|��{�{݄A�z��*ei@
�:���c�#;0���K�����U��7��#�c�t�:��%]����Q��M�9�g��{c���Q���c�{���Tw)�]�Y�u�f,µ�1�E���]�f�W��uM��7�9���y��n�Ecj��}�jGk�~��w���4$�Y�-3}=9P9���ő:D	b~^#�	��>	*RIA������}��?�ѾX��?�����A�� �������%!|���,� ����_���?�?AHs��L��CAFU�V����PK   㫦X`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   㫦X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   ��X���لO  �� /   images/cd9a76b9-8a14-4d7e-9261-140514b5ac3d.png�XS��7��*�QP��E�&EQz�Ì�( HWiCE:!0E���;�H�� !��)����y������޹������Y{����k�$�o�)m�rp�6嫗488��98�m���|��g���ʷ7�?�M���檎=��5�o�/p���p���➝	�}leno|��D���4�(w���0��n;GN�t�&w�M��?���\�^d�[ox�-�M�3Q��7�o�v��j���
'�S|�BjyI��00�m�5@/�$]{^�!��J�WW��o������3��~5�X����n�x�N�Xc�n�+���!�Y�[�ĩY|��/����(��NsHG/�ȤyxԆq�%�b2�R2vZ7�kR�u=�כV�Y�
;�����a=r��/�|ߑו�����Mkڃ?�o��.�Խ�;|���,����*���5B�ؖ7r&�E��nZz�������e��g��6}�bq���j�QRR2�k~[3�lM��Y��-,�_6m�h�q��U:?��v,
�H���1���&\��n�}�s�ti��]�vij^�	ٵ뵉ά�b1��D1繄���+z[�g����a�g�J�7_V�T��R3>��Y���qΉ�q�&0�������}wwy�H�]�j�ς�կ`�b�=73�c�yR�a�g����3�����~�τ�,J�f�hPt_�5�{ .������A������^�2���,+ϲ��k�i������N�p�ixy%�����XSl(���^"7/�������677���:.���;��������K.$RUS��ۚ9c���|�ϩD��K��n%v�OU��47��@'�3�A%���X	F�!�D�������(cOOE���}4��E�PQ�٦/z�#m`;C��r�*���Z�XP��*˄���OEbF�@ �.L��-�EJ��o�e.�c��JN��6��b�����~��+������l�&:��F��ͷ)���Z�?+���o�,�2-�/��Q����:Z�e7h>����Мf�����P�X|aH5�y~�J�����C�Ζ�jA���b��^ד�.����v�Ym�ȯlm�މ�M�(}UD�U�I��m��ͽS���>�����
�)bi�?"l���\&&&.�m�^#Ą�~7����S�P������2-�agC#��f���2q��I�ɡ��55oj���t�b<�p��f|��Ǟz:!�bO>�dp�z.]���YS���V_��\�c��X���#sY"����sCλ
Mu�Ė�|q��	�̗��(jX����d���m׹(��^4rj�#;'a�+�D��ͽ���2N���S��S�C4�JV���+ɹ͋{Щ}U����,ݾ��DA��"R	���k���2��Xn���N���;�:Ŷ�wBjy	�XE&`��[SP�rL��i��U�`7���7`�Mhpٕ�sY���P��l^y� �D�p|���Pfv���{VVm��L&�X6�h��}TKK����f�Sb���͡�H6Ťyqy�ciD��y�����n��׬�p�&�%�?I�Mf.4�z�ϒ���N�����(l�%Kd���������{�oii����TMg���y9��(�raH>��F��8�0�V5I׏�1��ك��}���C1�s:r��(.���Oc䅔U���g�X�]NUC�_�OG�_M�L�q�Ilz�דF0���w�g2�'��7^N?֞)����������!#��(A��]�y̺�,���o;te�O�|����(>&��v��q�W·q�F{w�{��B�?�4�=Ļ�e���fg���㭜��ǘË��[���®3f�޷+%�Ŕ3�Дv��w���գ��]tO*�:�aSa#YK`.v���U|�F�d��@9���y����kJ�H-���î�������\�if^���%W�ܗ��!����˃����w�C,U�.�7��/�4QI����dd�l��)��~���6�Ɋ,��4��$�2U�m����>2�Y��lf��t�iCtE�,bt���+�^��a�P��`�(���;���a
����0yF������j��>��f�����5����}�#���y��鱆ŀ�<k���<wi�:�v%99��LT�3a*��`�:�Ƥ-�q�x����?e%���-��`�Uh#���S���EEE��[YR�[��Տξ�˳�;���#���|�%V��X������D&�XU�4I{��:�8[�ܤqE�Kt��\���.��Š����/�,��a*��|�1��
-M��BG��������	op��CS�
������(���2��5bw����ğqB�G�P�f	3��%KӵaL�]v9[
prrb�j�����9!��?���$&ɣ��Z�����s�Y ���`{d���/�/�z^DEE�WgV�]��2�	+��}��������������Gnb�˞��)`�e�߉ZY'�5����m�W��Y�NnS�%{�����mF-���{�5��i@1���Ӹ�,���+ڃ�GVVV"�ԋ��K����,�)B#��=L9�S��A�6��v[�\s�<�:!�<�1���j��d�z+����/*T�[zr2H���}�Hi�2u���(���x��`�vS�.)4X"�2��
����v1��^gW�KK;���,%ŬY���u�M�7�џ=�\��]@�0�����g�H�؛��i�9x�~ȳfw��y�}���0���f���1t�B4+�r��|MBTZN.u�܏M�����`�07+0-{�6���YN�Dd�!)����	�e��A��A��p7ڞm{2�@����wt<�
����zbO�Ts�$�A���H���k���,�F�1*���{�x�[�u�o��6et}���O�rm?k"�����yK\�y)w��ň:ט�b���=L��l?g|`�50+�":������l�l��i)���p�؞�`����bf���VKz��w��~���KN�p�E��i�r��U�_��P{���,�D����9��gj�S@���vUv��}�8P1��<�h��]��80	�g��w�/1�e�M�
9���.{�"�����,�F<Ɣ�����'㒓ۻ�Tn��'�����dgE�66w^�x|brR�jąː�R`�6d�'�C��I�xiŔ����8���i4�b�AP�ϩ2�]س��O�dؼuH8���+,��,��L6�e���3�ˠ8�P� �vo��~�]S`.W�x�b#��]]IA���򗰨(>
3dK_���T���X��ʦG8k&�u+�6]��dP:�k��E:?9yx��V����ٷVTz�Viب�[#eU�UlR���F;�������ƥ�3�l�}V�Ŏ]QG$RSs-�L+�����D^+j���.��s�B�sخ�cW��3���tu?�{w�v����|�"cbl���M ��'�\.�ɺ�|e-+�}Yּ� I�|��nK@��6B�UֲU����ԏ9x��v�����Du�p�ɧ�1�{?� FI��y��/�ck촢��{AWX��_O�ð�\�=)hVΩ1�aǆ�8��j+��Jr[β���+%���^�	^^�m)�-��Ω2m*����GGo�]�2��wE�P���R��VMO]��`�j�{�#��!�׏��,��?A�6�1�O�#+���	ۚ��1���?���7����47ֱ=�ڲ�G����=�K�kV�\e���"��[�#0bl��e�}m�#.��Ҩ�*��A��4|w~�;�V�����Y�草͏��l��Odk���T�G�TV�@�Y�9F$���@�0,��N�H3o֮���I�6!&��(ё�}l����x`z ^�{y~$�bS�'�����ǿS�V)�/4�ܡ�?8�q������_�����ej��5e�q���Yu�!���L�Ql�\69�ᵍ�'�{�������f��:��0�-�NA��\O���x��0/t�.�f)w���j"QVb���@@a�f7�<g#��s%���s6$�b���셜}���Ma�H��"��'8��EVy��%Q�]�9h�r��FMx򨯟�_8��^��,����|��S��M�مOkY3�%�k�
u��/4���y`*٫�^6��6No���3Od��������:���'Ϩy�������h3���54T/��D�+���ND��qt^N��J����d����y]9Q�e�����Z'��--O�_�"[E�	��^��Z���
�raV�q*�� ��6�S�hY���l6�W`w���Ȫb���ۛ�x7���ҕ�N�����z���i>��^����L�������,Je|ݾ+���\3v�zy����5�	�]��9%�҂����.��d�nd��xKR�V�Yy��:�T�s,;�!��ʦ!KD��Z�J-1h�pE�=�,�i�W���,Q�d*�����LP��!��^�C��#�Y�Ȼ++d�,��:I�BL������6�W�<�h�t�4p��N���$P�����B�������%��qI�r4�{�b�M+b�W�q�S�V��g�Vb�r	JԠX��*����a�M�Y���f�%��	�ZY�����`w,
Ov=�Z�<N�*cc�es�☕Q��S�����ρ����g��\�z���\N�"�]��Q� ��m�pִ[�E��b����2ƾ�3��N���T��/�*Dy&ᾣ+��!F]��@>R�u0�޾:��Rk�is]箳頕F��H����d��N�弮��G:�B&'q�Q�iii�=û�o���W��"��Q�6Kd��1]������a�?���daGDD(�2�]���Gͼ.U����'���V:Ű�6K�����uL_�Z�^mq�H�}q�$�a���Y��[,�����'�}]J�ۧ��#��o3j���\��N�/�� O@����x��+�`��ҋD�S������^5���'@�_'���Sw� 8HA����4g�������{M!�$��(�V�hmְ=��xlc���W�����:�b@8c�Q�C�N����8w�Ձ�a��N�Q�U^�[zI)q(��2FG��(�q&�)f+���z��C�de�/wP���~PM�>׾bnn��Dg���EU�*�������'е}z��Wؓ�g��U�tt�a�L��7u�q��˛�Z;K{H��}@z�^�b2U�Q�R���Tɣ��Մt��?���sp���F��d0ga�vB�yy�6�u�ۘK�"�K�j��2#�fN�f[��^$�U���c�J�A�仒ǯw��F�m��>����Þ��?ZsW��Z�������������a�C��Q�NEG(�I�خ�z��E2�qb~^���V.��
 	V?��P�%Hד(-I�l';sV���уȑ%K���M�\&�j!��6�ȃC��jUU�����a�Q���EN��D"�n PR�$��O������^�	�h����~?��e�hr[n��U�)��|�#�hJ��=���-k��y��4�Xw�=ü�
�f\�$�f;4'��&��_$Y�>�8�>�@׼9i;=\�]�#�CmԤ���<#�X��1l�T(�D�.�C8����#��^�XQ�~�B��c�v�X!�o�����D�� ����F,�c���TJ�@�jVW�o�cQ�	`���N�1�!:�d���G��%E$4�?UVVfzH��_�MT��f� �f2�z�X+h�d��D�>���L+���W�͚�
`d�?�Ō9���N�l�ߧi�63/q~8H���зAG؃2��0V"���	���d�;�����
�Y�������K�hV�|mV��K"���_d̩h�Z8��o\ܣg0��QE���E����0|m��Ս��42���E�����+��ݰ�2L-f��6��ӽR�Fw�*�Y:H�������3W�r��84y�����ئ?%)*�;x��-�^�^�'ƈ�c��*8��ހ4:,"Ԋa�^;ۓk�w%4��bF��5ms��M�n�y��U�	]g�I�	y��f��5����4�|8��u�))1�.3:��Z��b���	3^.��
���H_�u��Ը�6��H��l�
�|��򣳺��K`3����"H�S#�w8���2��P��Z�!P T4���4=t�sw�1��0]�� A�M#�P��3ǈ������ޠ@M���"�b<ӳ���#;����;Rf�|���GR�?��],A�Br3�m����D��$�Kg��K%��7t'k�f���܊?�SKP%$��`��e�"E��Jqϱ,j�@'_Ŗ���n�F���Ά{�w ���9���O�����F��)�4��z��'����N�w�U�u���ʌlN��3_J`��{��D+�u���_.��Z�K��H39��ܒ(���B���d�B!�~�ub-B���"#˰$��@���,>����Nv7��p�NNs?}"Zv\�Tm�;�T�8���+jA��_�"�eF7ݦ.�@�A���GPn>˝����D455��D6�m͵tԧ�}�K�,�!�HGB[�
��������o
\�f�f�n���,��j'�J��5�fT0���������&IGy���'�0�6�j$���lOk'����uY�H���Ƣ��r-5[/5��~O=��I�y��xy�qWng.z�e#^ʼ72Ƽ�f�=�b
��d��ׯ��<������������}�}���o��6�ovQ���b�0Ϻ�?�i�W@�����`e%���۾}��ĄE�ъ
��q�i�L�"��r��$�Nq3�a�ё�8 m��BLCaz�^�U+I1��Mw�e��cO�}����ǂ��=��$3Ɉ4�TJ�����(Yį�L�O+�H�B�+��]����)��bZ�w>���I��q��ϊ��}������LX˃3I`�ł�����-y�_+�L��tC��js�+k7�Zy�P����*Ǚ��2rr��St���������sp��7Q�+�f�އu�I�;�&&&�Aj�l(B�P��#����_r��W<��k�v����[��� ��6D˧$�Ǵ55��@3�rPV�&u''&Z���W�3ؒ��򖓛{�8�ted�[���I3l[XXHVZR�	���֔saׁOn�!ӘaT��9��ٲ�x���RS�ua��<����4��vvUUU'}{�r����� !H]!	��B+�&����e�X�r

\�: 3>lu�2ڕ����N���KF�ZH"S��^������r�T�_nc��m��#�����eeS:,��,,긕�:�NǚSr-S���Wb�*p,Mg��֘�����V�F�V��d��1^?�ztf�c��V=�s�#8��������@x <����@x <�} �*��y��u:/��p���N�gz`#�F�N4�Jݶ�,�_I/�F0��`#�F0���g���OF�[���U�*�z�#�F0��`#�F0��`#��G���W��+��F&:3���'���q����_�#�F0��`#�F0��`#�m�}��*Ϧ_oR�y��uod*�o�������V�Oi
��i���>��j�/�^�A��?���c��W����U��a��@X ,��a�m�v��K+������a��@X���yy��r��������8�0^�g����X;R]��C%�"�+�����'��G�J^+��Dj����'�=ڹ����N=��WS9~���ШqᲺ��W??�ͱ�܍��A��j��瘇S�NY�]<ߌ�W��?Ç�.rK�rt��\76N(���ҊE�C���RE=n�3��Y�С�!�Gq1ٕ6������P�TDm�UR�B<��|b�������bm��W�Kt��Ε�{��?vX$<Ohnn.3�8<���9��T�hLD>��a벯^���!�C���ώ��I;��ȗ�k�ߙ�$�XI�r~�%�$,�kr���2X�O4r����	n���%�,�k�!�g��C�������a��@X ,����lfٗV�`#3�$62���ӯ0w��+b�[=0�,Fb&�\!�8���s�_�1ەv�=�N}��b2!�I�9GN�#K�O@߿w�Ǻ�◽J�=�V˺����M�L�w���+PC�V�a�T��s�CN=&�w�����:9�I�)�0d$��4����:wb���Vzv3��g��Le�����Z�PDQj�p6�0T��Ɓ����`�b�
L1G���	��+(�]�L��']���T�sP{�0��� �ǻW}�����,�w�U�ȩ���{���w�?<�}��ѭ��	
/��P�l���uO�������?�����9�:d�v�IߠN����@X ,���@rҋ��g���a��@X ,�'�-���B����$i9J~]��(&�'�>z�W�ڬ�h�uV[�`�2O�jh�zj���W��yG�ʝ�)��_U<���e�"1R��"�8��F�,{�,M/���sj'{P��Kxj�u������v.s۽��.��C2M�B��E��T�ù�����l�F3�2�V	l'E��-Z`�	9޴�YiO���À�%��=�(�F�(����Z�b�C)b;�v~S6�Rҧ�ɜ@6�>_���?������z�~���,��/{�@X ,��a�����",�n�\�9�-w����oD�|��ݛ�З�y�����.�c��x��V�a���� ��`7O���.�[z+�M�׾O�H�5ڻ��~�Z���r��+��r	���r�������o�wp8[bh��z�i�wv��*/bES/�9����'н_��fc/:�㻛J�x����;N,�����6t����)iF����@�QKl�8���2@;�D�r��Yh�+G����x��~��)�ӫ����X ,���7:�ĻC���
��a������_����-�`#�F0��`#�F0��`�c�70.9�ԍ�l������[�F0��`��&Jx�i	}௢�`#�F0�����O�|\��N�EW�nb\���F0��`#�F0��`#�F0���N�ڌk�W�Y��J�nf�~�F0�[#��کU���F0��`#�F0��`#�+х�R2�e��2��`#�F0��`#�F�A��fH�Y���^0����_A��&�wR�F0��`#�F0��`#�����KɌ~��`&�`#�F0��������m���E��`#�F0�ۢ��ʸ~��N
#�F0��`#�F0��`#�}Q�y�Zƥ�RZbf����7�wv���`�?��-]V=��F0��`#�F0��`#}G�qj��۩��zt�MP>i��Yڃ��#*q��յ/�x�4#�~�/g�f	�%Y�W���3��s�`b�`���G�2?����L�������������!7c6Z/װ��2V�x����&�:�~)�~]|��u�z+?�:c���L�0����j��a�s�gjۺ���;�?�`@�@�IO�W�E���7�	������6��عť�Ԓ��8�Ϣ54�M�cS��:)������r�{��!)��p��y�76ځ�$�h�Թ-^M��j���*�W���7���������kybJ<۾�+Xz�I,��c�v�-�����5������y�8rG뭠�]V����Fn	K���7
{k����� +���f	���o7���ܑԹ�k*|O~��:95�o�B|Zåޞ�G��hqe;�&7��q8E�����޲�ߪ�����j���c�p���r���U����"�

��8	z�e5y���b��7�R���������o�ȅ���`���dZ����y�7'������by-��@F*�<��P��
���\+�[ȵ��C�л� �ˊBu�7��;�b�Na�Ah]kX+��o�"۶S����?8�\�L5�Dr~cP����H��P��N`��	`���i�s�7��S�}��ޛ�am�� �]�>1S%�m�$�ڋ�ϭ�����zt��z�|�����[P�Ruν�uJK�_�����7��c��^�f����W���h��y␹XǑ�΋^2�N�mP��1N*��/��B�s�	�]Y	s[�Q]��+��r��2F[�ۀ��8��	!Ae�bs�JUߟ\�aؿ}�Da���dg��b���1�^����m}�!,���u��lǚq<�մX�7��'F��1�\*:L��|�cS���k�]p]�&��x(��|Xk�g~L��s�̠5��7@��0렘Wl�q������_�ud������'��ˡ�a��^�V�V�V��)����fA���T�0^����P�sUd�"���Vk�}m2���呺+Z�y�/sآ���
��O�x^�*�,e�E���^�q P��{"�JЅ·��mF}r�}Vb(����k�LE-IQs�'.\lK��FZ��A4=�M%�G8�'��2�f����wQ)��Bzo�9��6���u��ha�$C�����Rt��Ķ�p
i(yWf��m)�e�	�٣�'z��*���ߝϖ�-�����:`��~q�YX����:�NW"8�{��c�=�[�9�kZ�FQo]K����R����ʴE��¹��~�0dw̦Ϟ�>�~gcB��:��	H�2!�o���N�5�첢��b�p�G��g���C��C��ЕA�g��u͘[c߯��^=��xBM�i�f�e�_9=G�m���������˃t�vR��<Ց�%�C�[�H���.z�2y��"{��		�6�k 77f�/�h�8�����N�:��<UB����ܞ<�m��	�)��i�t�c<�<�,fmÝ������.�hz�\�<�[���}<����י��2��R�ב��;3����R�%��s����o6]8#�Ӏ�+��q�%#u�4m<�	rQ8��-�m���+*-z3~4\�V]�5k�6�݇m���y
&���`x]]�[��	,:�p�p�V�`�����!)�"�p�t_���_N�7�oT3�ϐVK vV�t!N=�yh,=���zب#"j'�`sYa>�F�F��ҷu��3������ƥx�'�n�h	*��'�^�o˰붙�m/R0\XT�
�C0WC���U�h����@�[��K��D:����(ؐj��_"vddF�-��Yh*��i���5`ĵ���s���F�wc���5�p�n{�J�z��F�t���Z]������r���'��+�F���k�@9��j��h�)�q�G�/����k?D�7�@��X�*����-a6�Ԁ�y`p��o�����uWHDo��D3���k_B�t�9Ɠ���&�m]�=h������3��8����_o��)�D��f.�qyr�e���3�#[L�B�(���ي�i}.�=���)�8��C��-Ϳ
�=��%;������t��o�ܲ�}���^�f��y��DҖ�����@y���缓�����X�0���ȶ��H����H��w�:�\��.*���/~3;#R?��X(I?����=�qX�����R�|Y�ZJ�� ��]饌%���i}1�=�e����rsþ.Ϲgf3Cg�Q<5�u6gf�BRi���ͳu��#$S����Я��^�������8s�)n�K�rJfD�`�;�t7����oA.��.on��|�GJ���x���շ���VT��8���1ZYf����ڬ㉷hCET/�����o|H�$ta��#�7t6��hC�$��;��ť�4
���y����b������z���û\�w�� ��a�O,�LY@�83Z��v��=��v�?4fg��帞@<A���]4\���\�4�Rt��+�A�4��%e��|u���/{ژ<���),\
L�R���=/��O�]��SH�� A�>�^��c�]��*�G�+���<U.Ut���é����[�`��'Ԗ�Vψ�٫��[��쒥�p���Q�H󱡁K��w�4�K���h�t�h	���Z��9W��d����'���9!/o8���{�'Ч��m���#p��u4��������Z�P�fh A��~dxH��;U�Q?�*�*wB��Q�������<�~yB5��uS�ξ��Q�RA����\��PQ��P;�F�>��cP/�S��w���qo�n��܍��/��'v܆D��
�������V2&���ލ�����}ת�U���^��ܪ�ڗkKw���:B�$�*���wb�E�c�=��e�z�*g+���������Z�Z���sV��%*:zy�gO��'����\��˪����N��[r�k;-��n�� ��҆��n�V�n^u ��*�	�>H����gl>}�^���w��|
=�5�P���t��������K啯!l�>A�Bܥ�ң�	5),	�A�pwV�1*�NW(84}3�����>U�+Kt��/P8��_Ҝ�z�hχ����z�� 7R��g*K�q���G��|]�Cx�|�辨��bc+�O�������@;�C�m��� 6Zx+k�yd6@���ّv9o�w{7��s)G0@t�2�Nd̤��������~��;
E�N�@��ᾦ�׎���V.�jҪ���oVpٗ�3Y�>E�#���a�F/4ħ�]����Ju�F��y#&:����v�8aKMAi����
����M�-]T�+aȲ���Z�{!a^z�V� Qa��y�b�P����T�)�	THlo�����}��e7*!72�f]�Ŷ�ȗ;WG{S�����sA�?�R�7����C:x�ߣ�vэ �煥�޳K�o�zF�j�Bn>2���/w�h\K�ߨ�<�D���a����I�Cz�I��v
$����>����K_��m蚾d�賠��0124�R�6pc%E���VM̎�(���8ꄦ@���[���'�@�C���h�x<%��׸����C�h�����?����_��X�1�Ȩ�_�]�� S���!U	��Rt��ρC��R����ȅ&��<�B+@l�������%A�������1�.{Q��@K�^���x�KK�6NO�dD�����B��W�:��
�Y��x���z5� �I�f��~�k���ۺ��竹b� w�2�mf�����JX��p���S��]>`�"�õ
C�8���y|M����kJtf���Ly����F����'<ύ�C(x¨yB�����_�@wT�B�G��X�R�m��Z0�Tĉ�q�zh	s�VH/��"K$��+w3�qi�}��Q��GwM�N��9~�T:B�Ae��$ϊ����x��Zuϐ4.��kB��Ӈ*��W�4�(�L�n��F7���S|1<�'�ۺQ����WW�@�-n�CO�(��-\�2�͈�昫�_� �cTfppv&�V@f�Խ�R�]Rab5ŽBј��6u�C���Aq}�e�j7�lȲ �Z�������K�ڐ�@�V�C�f�=?��D�3������� ���O��������2Z������W����+�E0�5K�
l>��W�aK-�V��l0@��	583+�ae���O�z��fM�OB�I��� !i_�cuR�r?Ŝ�;>I΁��T�	m3�i���R����9��'����^�PX
�Fk�Ʈ-xw�B	�6���15#A��=+T@��,��ǽ+���YO���h�s�U�b<�d �V�N��P4�X��[��5�DOnT�{0y����	���x����
�%�9���yB��^K�g�od�vi��	;���C?�`���2-w��W7�.�9b��4�x��io��շ<鈼����';���Mi��9�O�K�©y;.auwڽ]���(S��go��g�h��'��#��#~iGK�9����wT:Z
���5?�O=�$�����`�9��ݱ�晻#v,zFW�U��[K=���qӷ�F�M V��sH=�1R7�C�3�p�F�K�z�َ!�d��Xo~��-ѝ*zP�o�0�<g�;a�ck(s��f�I������5��}��m%1�QK��2!$��OT���t��4�P�?�6����fS�:P����X��ANtac��X�A㍳�T�o�'³�_�Pc�ݚ��hIm�E�;9�x�tb$=��oG���@>�Wez5ٺ�a-zMLn��8��~5����P*� S�{�k�]��F�ÜD�,�Ʉ	�֫�^h�U�����!:gp>K�ʕQ���U_���"����.��p�h��	\t4V�J|�|�Rh칕5cDl��*'�Lp�;�r���I��e�=���ʖ=����SN�k�x��1_��
�R)V,W�j�T������.l����e�-Vi�~��,ntԠm�(�e��չ�`��|�|�:%����Z����7�l�@ݚ�_��nr���������tw7ƒ(D�5��jn҂��u)4ѹ��(J��i=�h&[Bӣ���/�5u7�n�I�3@d/��A7�\I�tϗ��54��xS�`�#���^�^	�OӃ�o$|�������NZԂ���;GhA�#	u0�{��m�OM#؈>IA�L?_����7�+��.|��uѲ��O�zRW�Ȫ	Ww��v+�T�-> ����wQ���T���B�r�A�V,�-tGW���?@V�T�	��@)���z1����v`������d��t���5T��Xpל���4���`�3���P��*y���r��d���B߃N��}8�<-�j"�?�|RX��Ox�p���c秿f�ǭ��_������N�=�����S�Ni����^5E����܇�=iG��������2M`��9-U��� )�1����� �Hz�Ҙ)[�����U
�O?�]G�HX�MP���YA���h$�� �N�m�c5�NPG�e�_��kU~Ƚ�B�<�fn��j+#0��隁��4#���������2rMV�R,}N�#Ա�y�m�%K�m�N��I붛\4�ԓB�:B��Rt���=zy�s�r�N����2�j�pw
�_�ײ�fk�|��EAt�ʸ��kdW���=*gs�_��zӶF_I~*��Ze���{W��0\N�#˛�6���"�������3��ٶ}�F����.�٬a\Pwo!�OҾM|K��0V��8��ݤ���Kb���*_V���GR�,q/���e��ef7�sbdǪ *G�\O�qQ'���������[�vB�<3�A�ӂ�����*�I2aE\P.i�j�s-�/ۼzF%l<o;>��̻��?T�����u� R/�y�US�1�?���PiΌ�]bX+�ݳ��"$�"��| �S E8�v.Q�vҰI��,U�Ts�;Ϭ�l�0�k����s]�pdf���uT�c�c�v[��0AªY�N(~<�i�KWk�Z�n���I��7-�UՀSI�W6׼�@�,�o\D�@�Ɇ�f�E���1�	p�S]v��E;�g�Է�����]��y�i���*Y�Рl��>�@�=��k��;+c�țg�la�l�\|�Z�>�~�'ե��<9��*�%��܁�D+)υ|A�%�4�[
Mv�x��4�h�

5Ĝ���x�xx^�d�ﱳ�����f����:���7A͞�2Ư ���같��Bh�nT;� pR8���и�A����C�Ñ��Q�Gr|$��mq�������3�	.�O��%�f���!'Y��"(����r,�8.�X1?���E���-����H����R��{lz(�K�6
Mc/2�$B�J�
0|����ЎX�Ƣq��*��1�n����y&�X�q"m��ֹ4S��swuo�=�������˼���f\o������z��}�Pe����Û
�z��9��W!�L�J曚<�{�鯆?����c&�B���r��4��aO�k���(�m��Q�UZS'��84x�f%���t?�����z�����໫R���Y�Ң�lR�$W�ʆ�7������^��rt'�r~�l�}����h����v�D<�X�p$ۃ�G�.�B�؆~m:ZWɳ-��ށ|��*ywW
��d�E�`�] ��}=�J.m��lP"��<��I��l[��^���r�Hp�{���G�Q�����8�.(�O��q*p����`� +�ԭ݇R&�w��(��i}�N��kʖQYoɺE����U��&��*���\zj���_vuٗ�/:Y��g/�C�NJ�='84�`��P�n�?8V�Yuٸ��)g�A�ۚ�.D~��<L*g� ]􎯫~)�eZK���O��QK� {Cs���'���J���B#��Y]H�)Pۭ�q�ʑ�bINP���D�ZZqKŏW'�t���-q �nK���OW�o��B���F�F���M�Ƙ���Y�g_3j�����j��A]�.�E��|!�@me"�W�7�������܁<�χ�* 	��f�������2�n�*u/��h9���f�lw	�$c=�تcRh���O���d	�k�%��Xh�_��3K�<$�2Z�v�]���n<��~i �(����������3|���2!g{i����X�54z�P��;F�ɳ�J���ە�����)�������cUT���*C���<<�#�P_������,Ǵ,]�ڤ}�P,'ZR��6�3'��jY�+=�X��`�������Z,_'���g@���A7�N_~�Y���$7(�˹��Rml�ܯ~fĜ�d냏И����X�f�ʜ����
��:�;Q��vP-��[��1��.��B�9_��=Y���^P`
���?%-<
;�cܭн�ۧ{���'{���w2��9kA�/g:rw��� v6�,�t�������u'���t%�iz�<�D�:s,*��2�����c�k�ph�~�i�	�u�˿�Ga-�Sڊ���A�?��?'�2�>�a�3y��<�ɝI&��S\�U��E���Ӗޙ;j�9��,gu76ֿ��3T�y���AF>c�)L�臭��"
*?D�Χ�/
+�7Aʫ"VѦ[�}�<�����4��n;��j�N		_r�N�SCet��+&,�	m����ү���Eu��Isq�O��t趨��Nn��@��/���@]�K����H�����k�f�'�M�c�!n��4��]�J�v�Qr��W"WM�zmkn�pbAl�i+�r~��Β��*���T��fO�I4w*O̲aw��Ҩ����p�)����Z���x=������X����ҙ�g�ϴZ�]���6�*�+o�3�.n��F}!��+�<z�2�4=^N"靖\+g�a�v���	ѭ������w��]U�nn�d�|��ׯJ�nSޡ5�C&t���p��~�H#��Q!
@k݅=R�Ғ
�������k������.��s���&�����"=��.�m@lO��w���hQZ\�*�a�q0.���#.��;�[6�w�%��@٣��>-8sT�sk'^E�G��5m��I�1��=*��B`�L!�G���i���_W��h�)�Z�����T>/Q}� 9,�S��M�
9�T��t��Ab�gk��Mᯥ��CWg#!�t�Ϧ�)_����*�J�6���5��D^󇖴R�Ns���j|����l�9ۍ�tΟ����0.?+/��<b!��}Sd��"Ё�v�q��7��b#Rg�b*㕂JP/k���#B��<���Ⲳ�+4�W�X�ZK�uQ��������9���!�a���3�\�5�2&U9-���'0o�3�,�]I�Y�|��l��*|��-�l�YdkX�x���i�r�G�F<�i���})�Rtϼ'ѡs�m==Џ��\E�A_h=�A�E��t�Ji�mLO���1�'���F���V����𬰮O��{��3Ⱦ�:zFS%�����=�4��Bٝ����J�����p݅�G�򵎷�܂�?@\~Ai")gi䪘���n��i�F��%K�Z���tb\4��Q�xu�9râ#��",��T�q{�ً!�XE��]h\[x��� ԕ\�O5�~"=+�s`�R8n�Y�xz-���2O�h����1]��uA�-���Ȏ�����3����7���z��Mi�;�*���o-]��ˈ����[�����[�좼ݺ��~6#��\�um�WZ2sA� J�#���Dťg�*�Ɓ���W� ��L�Z7�it��t�N����c���rR�����Z'\��Ljk��k��?Kؘ�,r���T�U�ڻ��U]�֣����3�4�w��!���r��H�Wû s���B֝�Fk�q�9����ڻ��$�8N�Z�i��͝�nJ��y�H��6D:Xt��$���LG�h�m]�mI=(z�`M�,^�B)w�3�R�����0i� f��%�������v����=�����������}� m���Y��ŏ\�Gֆ�e�E�j*�4���I[e�����B�g�|�}���<�0\����ߥ��R�"���i�X;Y'���Q!V�tܼ�'Eq�ڸ�bx����t�;��v�?���H�4�������M�p �������ܕ*�V.�ʩ���J/z�י/1�S�������.��5�2��F19����<2�o]��*��S�ǆ`X�o=��Hd�܍ELV~b��7U5ͽM��9
!��Y�����VM����=ZR[�R�5��\_Q�Ύ�������"�����(I-�oE�G�.E���6��6�I��ȁ�Z��B�!S��)��n0!��=��#�5DL��>�o��%ĨϸG�h]�.L&(�Z⛕c_�UZw+�6d�DΝ5��@����G��đoj�@J�/Dm��+:���o1Z rE��LqZ��Y��G�[U� -Ab\�+�f�T�GK�����l�9b��
�%����4�n'6�*�%�Ax�Q�Q�4��N��w�q���V˾yf�Ynfg���+]��r��g�f�wۚ7��#X"%m2�jk���I�B�>ss[vr<gKO�.O���7	f���ToK[W���N	����&� ��sˌX��G\�T�m�ǵ 9 Oy��<�9a��$nS��Y&�>�X7};>�NȪx�����"��I`��%;m*1�-���D:M-{������Ъ�,����6Ǟ�NޟZ&5��1,�;n���/M?p��`NwqCQ�e�����R�ZFJ�8o�m�xYTϧ��3��4���S��1	���N���CC���=2	0 ��,K�
�6�9���O?R���z�x��E2���������PX� kY��w��RCxL[�P��ܥ������"e���ke11M�v���t���SP\pު�N��=��A�1�ʘ�jsd�^5�{�o;��9%g���^핯l�i�%�|�;8���]�d�h�_�N s�bC�Vn��(I���LbG#���{x=U?3"�t_iOm�ԧ��G(�y=�B�﵍R��v�u���	�&�R�^.FV����������ib�쯬����j�SS����q�c@�R�u�h��B�>Wj�"ҽ�>���9�X�|d����{J��] D6Z��Ƿشם�L�P���-~�	D���0B���3\xc���ɴd!�D�������Q��U�z !AB�� !AB���iԷ���T=W���� ����!B��k��;r�w
-��M�I��;>ߋ��Ye�,J���.�ݳs��܄��V�Z��G���'������C͂B!��E�ԪG�`���ιL�<�s� 'ՓI?v�&�b�"N&��Ѱr��(��%��^4W����*خ���`m3+��e�ë�8Mje�Ū�8�scl�Ӳ �ˌ:z�rȋ]l�}�@��('�<�5�H�;,���nl�D����XT��K�*؟�纳�Lc�`�l�l�\ _��m�e����9ѓ�o.��KްMeMs��,��t0���y�86���`�VLq�}��|_P״5�p���>$| �L��PK   㫦X~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   㫦X�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   㫦XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ��X-�T��  
$     jsons/user_defined.json�Z]o�6�+�_g
��țWwC�&)�&/C0P$�
p$W�E���dgY#Q����9u�u��9d���ϛ0?�ﶡ�͇����/�B�-�
n�g�lwy7t;?�������{v��]Yճ��+�l���g8�(]S��j�z���~�Z�v��y	?��\p̐#űC���%��9�Uغ�ܴ�$���-�]p�51����WH� ��T8��M��+>��ݿÙ�Ԝ�nl��*��ٗy�{X����~~U��]�&0���u��_'�����ʏ;Ȩ:�7mSB8��n@�-��/�5\!L��ݍr��܇��G�gm���Y�<t�n/oo^��_�d��aS��{~u���(,$��m�ae,��]�QU��c�!�N���2�����mP5 �8	���@��&�.q�1#x�I��?�M��%��IEӪ��CJѴ�_�8�P4���":�1xA�QЛWo�#���ev�S$v9� ɐV���N���EX�Lא[���Ɖ@G-�
'-Y�d*l��БEK%8�Ț�Quuȱ�k���8�c�$��8�b�b���2td�b���HG.���Y�D"j�]ld풉�qr���K%���{�n����Wx
��^`;�$׌"�G���L���Z�<c�A`o�z��<X����������v��d�eWp�n�A����W��揌;/qWn�|��ք��>�^@w��h�]a]�k���)����a<RW�j���Y|��Û|�޼����7g݇��o͕���h�6����[���8*��@s�����H3��ŕKuT�)���Hs���9 � -�
{y���U"$��r��+$�[��X!Gce!rb�*�p[�e�M�W��s�T�EuF�"dA�� ���1a��)��O�׸_C���C�x�C� �W�m���vv^�]�$�_!�M�U]�T�ڵ�];ɥ<�s�|�CP/HXUP/fJ�r�yc��Җ@��* C%��cAx.�c~H���mmӾ}��u&��d����v�B�c�!<�Z�jz��ʄO�A/(�RyO�g ��f�6d���3�Dd�r��=ԟlW��o�wa��=�q��1�zd	����K0�%e�3{���������s�5�r�z5{�ۺ����Կ���U>8+�BB�6��x�e�_:(�X(L*a��s��G�k�(0ʽĈc^xku!�b P=$)*��`cG�"
Y('e�@�����2~�w�@5����,�ؐ#GW����X�U�1�b���#�3�3���`
(7G�	���w_'��T�����6����b<��C�d�6b�ˈ���������s���k�oe��Qn����6P@�+%F���C�/�藋����#�$�!�}Mb���!�є����(�X� �/'K�!�� 'S�_,��1?�<a�N9� x?U R#�_N����*9D`'D�����A����	&��GX���ڨ"L�����ҿ���.�����7T���:����������6aF3<��m�:�nB��_
�[Hh����RH2\м�*�C�y�A8�E`6�ݾ�W{M�$�@�{�D��L:8d�eH�� �YC�P2�<�&�`�8�����9@2M����#��g�|���މ�J
�Q���+`I�숢�;�<AP)�;E�E�I2l��{sfK�}y������_PK
   ��X)$�  �                   cirkitFile.jsonPK
   
��X[�o��� �� /               images/055d5e06-61e9-48ec-9da3-6ebf1aca914f.pngPK
   ��X����	  P  /             � images/471995ad-a105-47c5-9945-45370623043a.pngPK
   㫦X����+  J  /             � images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   
��X���Ʊ N� /             �� images/8eec4e94-481e-4d4e-9432-645515506382.pngPK
   㫦X`$} [ /             �h images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK
   㫦X$7h�!  �!  /             � images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   ��X���لO  �� /             J images/cd9a76b9-8a14-4d7e-9261-140514b5ac3d.pngPK
   㫦X~��a� ٮ /             X images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   㫦X�+�s;  z;  /             � images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK
   㫦XP��/�  ǽ  /             �H images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ��X-�T��  
$               �� jsons/user_defined.jsonPK      $  �   